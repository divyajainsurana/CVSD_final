`timescale 1ns/10ps
`define SDFFILE     "./MEMC_syn.sdf"        // Modify your sdf file name
`define PAT1        "../Patterns/pattern_MrPickles_gray_4s_sr5.hex"
`define PAT1_1      "../Patterns/pattern_MrPickles_gray_4s_sr5_flip1.hex"
`define PAT1_2      "../Patterns/pattern_MrPickles_gray_4s_sr5_flip2.hex"
`define PAT2        "../Patterns/pattern_RickandMorty_gray_2s_sr5.hex"
`define PAT2_0      "../Patterns/pattern_RickandMorty_gray_2s_sr5_flip0.hex"
`define PAT2_1      "../Patterns/pattern_RickandMorty_gray_2s_sr5_flip1.hex"
`define PAT2_2      "../Patterns/pattern_RickandMorty_gray_2s_sr5_flip2.hex"
`define PERIOD  4                          // You can modify the clock period to improve the design performance
`define TEST_FRAME_AMOUNT 10
`define FRAME_M 48
`define FRAME_N 64
`define BLOCK_SIZE 8
`define SEARCH_RANGE 7 // +7 ~ -7
`define PSNR_BASELINE 23
`define MAX_LATENCY 100000000



module tb;
    // input
    reg clk;
    reg rst_n;
    reg pixel_valid;
    reg [7:0] pixel;
    // otuput
    wire busy;
    wire mv_valid;
    wire [7:0] mv;
    wire [5:0] mv_addr;

    // memory
    reg [7:0]   pat_mem[0:`FRAME_M*`FRAME_N*`TEST_FRAME_AMOUNT-1]; // 48*64*10
    reg signed [3:0] mv_i, mv_j;
    reg [7:0] mv_mem[0:(`FRAME_M/`BLOCK_SIZE)-1][0:(`FRAME_N/`BLOCK_SIZE)-1];

    integer i,j,k,l;
    integer pixel_count;
    integer pat_frame_count;
    integer ans_frame_count;
    integer block_i, block_j;
    integer mv_count;
    integer latency_period_count;

    integer pat_video[0:`TEST_FRAME_AMOUNT-1][0:`FRAME_M*`FRAME_N-1]; // 10*3072
    integer ref1_frame_padded[0:`FRAME_M+`SEARCH_RANGE*2-1][0:`FRAME_N+`SEARCH_RANGE*2-1];
    integer compressed1_frame_padded[0:`FRAME_M+`SEARCH_RANGE*2-1][0:`FRAME_N+`SEARCH_RANGE*2-1];
    integer compressed_frame[0:`FRAME_M-1][0:`FRAME_N-1];

    real PSNR_per_frame;
    real PSNR_total;

    integer SAD_per_frame;
    integer SAD_total;


    wire [31:0] debug_pixel_count = pixel_count;


    MEMC u_MEMC(
        .clk            (clk),
        .rst_n          (rst_n),
        .pixel_valid    (pixel_valid),
        .pixel          (pixel),
        .busy           (busy),
        .mv_valid       (mv_valid),
        .mv             (mv),
        .mv_addr        (mv_addr)
    );

    `ifdef SDF
       initial $sdf_annotate(`SDFFILE, u_MEMC );
    `endif

    initial begin // mem initialization
        `ifdef TB2
            $readmemh (`PAT2, pat_mem);
        `elsif TB2_1
            $readmemh (`PAT2_1, pat_mem);
        `elsif TB2_2
            $readmemh (`PAT2_2, pat_mem);
        `elsif TB2_0
            $readmemh (`PAT2_0, pat_mem);
        `elsif TB1_1
            $readmemh (`PAT1_1, pat_mem);
        `elsif TB1_2
            $readmemh (`PAT1_2, pat_mem);
        `else
            $readmemh (`PAT1, pat_mem);
        `endif


        for (i=0;i<`TEST_FRAME_AMOUNT;i=i+1) begin
            for (j=0;j<`FRAME_M*`FRAME_N;j=j+1) begin
                pat_video[i][j] = pat_mem[i*`FRAME_M*`FRAME_N+j];
            end
        end

        for (i=0;i<`FRAME_M/`BLOCK_SIZE;i=i+1) begin
            for (j=0;j<`FRAME_N/`BLOCK_SIZE;j=j+1) begin
                mv_mem[i][j] = 8'dx;
            end
        end
    end

    initial begin
        $fsdbDumpfile("MEMC.fsdb");
        $fsdbDumpvars;
        $fsdbDumpMDA;
    end

    initial begin
        clk = 0;
        rst_n = 1;
        pixel_valid = 0;
        pixel = 0;
        pixel_count = 0;
        pat_frame_count = 0;
        ans_frame_count = 0;
        block_i = 0;
        block_j = 0;
        mv_count = 0;
        SAD_per_frame = 0;
        SAD_total = 0;


        // output answer check
        for (i=0;i<`FRAME_M+`SEARCH_RANGE*2;i=i+1) begin
            for (j=0;j<`FRAME_N+`SEARCH_RANGE*2;j=j+1) begin
                compressed1_frame_padded[i][j] = 0;
            end
        end
        for (i=0;i<`FRAME_M;i=i+1) begin
            for (j=0;j<`FRAME_N;j=j+1) begin
                compressed1_frame_padded[`SEARCH_RANGE + i][`SEARCH_RANGE + j] = pat_video[0][i*`FRAME_N + j];
            end
        end
    end


    always begin #(`PERIOD/2) clk = ~clk; end



    // input state
    initial begin
        $display("-----------------------------------------------------\n");
        $display("START!!! Simulation Start .....\n");
        $display("-----------------------------------------------------\n");
        #7 rst_n = 0;
        #`PERIOD rst_n = 1;
        repeat(2)@(negedge clk);
        
        
        while(1) begin
            @(negedge clk);
            if (pixel_count == `TEST_FRAME_AMOUNT*3072) begin
                pixel_valid = 0;
            end
            else begin
                pixel_valid = 1;
                pixel = pat_mem[pixel_count];
                if (busy==0) begin
                    pixel_count = pixel_count + 1;
                    if (pixel_count%3072==0) begin
                        $display("--------------------- frame %0d input success ---------------------\n", pat_frame_count + 1);
                        pat_frame_count = pat_frame_count + 1;
                    end
                end
            end
        end
    end


    integer temp_pixel;
    integer temp_abs;
    //output state
    initial begin

        @(negedge rst_n);

        while(1) begin
            @(negedge clk);
            if (mv_valid) begin

                if (|mv === 1'dx || |mv_addr === 1'dx) begin
                    $display("================ Failed... Encounter unknown output data!!! Your mv_addr = %d, mv = %d ================\n", mv_addr, mv);
                    you_failed_image;
                    $finish;
                end

                block_i = mv_addr[5-:3];
                block_j = mv_addr[2-:3];
                mv_mem[block_i][block_j] = mv;
                // {mv_i, mv_j} = mv;
                // for (k=0;k<`BLOCK_SIZE;k=k+1) begin
                //     for (l=0;l<`BLOCK_SIZE;l=l+1) begin

                //         temp_pixel = compressed1_frame_padded[`SEARCH_RANGE + block_i*`BLOCK_SIZE + $signed(mv_i) + k][`SEARCH_RANGE + block_j*`BLOCK_SIZE + $signed(mv_j) + l];
                //         compressed_frame[block_i*`BLOCK_SIZE + k][block_j*`BLOCK_SIZE + l] = temp_pixel;
                //         temp_abs = $abs(temp_pixel - pat_video[ans_frame_count+1][(block_i*`BLOCK_SIZE + k)*`FRAME_N + (block_j*`BLOCK_SIZE + l)]);
                //         SAD_per_frame = SAD_per_frame + temp_abs*temp_abs;
                //         SAD_total = SAD_total + temp_abs*temp_abs;
                //     end
                // end
                mv_count = mv_count + 1;



                if (mv_count%48==0) begin // 1 frame motion vectors
                    // $display("mv_count = %d",mv_count);
                    mv_count = 0;

                    ans_frame_count = ans_frame_count + 1;
                    $display("ans_frame_count = %d",ans_frame_count);

                    // v3 updated begin
                    for (i=0;i<`FRAME_M/`BLOCK_SIZE;i=i+1) begin
                        for (j=0;j<`FRAME_N/`BLOCK_SIZE;j=j+1) begin
                            
                            if (|mv_mem[i][j] === 1'dx) begin // unknown check
                                $display("================ Failed... Encounter unknown output data!!! Your mv_addr = %d, mv = %d ================\n", mv_addr, mv);
                                you_failed_image;
                                $finish;
                            end
                            {mv_i, mv_j} = mv_mem[i][j];
                            // $display("mv_i = %d, mv_j = %d", $signed(mv_i), $signed(mv_j));
                            mv_mem[i][j] = 8'dx;

                            
                            for (k=0;k<`BLOCK_SIZE;k=k+1) begin
                                for (l=0;l<`BLOCK_SIZE;l=l+1) begin

                                    temp_pixel = compressed1_frame_padded[`SEARCH_RANGE + i*`BLOCK_SIZE + $signed(mv_i) + k][`SEARCH_RANGE + j*`BLOCK_SIZE + $signed(mv_j) + l];
                                    compressed_frame[i*`BLOCK_SIZE + k][j*`BLOCK_SIZE + l] = temp_pixel;
                                    temp_abs = $abs(temp_pixel - pat_video[ans_frame_count][(i*`BLOCK_SIZE + k)*`FRAME_N + (j*`BLOCK_SIZE + l)]);
                                    SAD_per_frame = SAD_per_frame + temp_abs*temp_abs;
                                    SAD_total = SAD_total + temp_abs*temp_abs;
                                end
                            end
                        end
                    end

                    // v3 updated end



                    for (i=0;i<`FRAME_M;i=i+1) begin
                        for (j=0;j<`FRAME_N;j=j+1) begin
                            compressed1_frame_padded[i+`SEARCH_RANGE][j+`SEARCH_RANGE] = compressed_frame[i][j];
                        end
                    end

                    PSNR_per_frame = 10*$log10((255.0**2)/($itor(SAD_per_frame)/3072.0));
                    $display("..................... PSNR of frame %0d = %f, SAD_per_frame = %0d \n", ans_frame_count, PSNR_per_frame, SAD_per_frame);
                    SAD_per_frame = 0;

                    if (ans_frame_count==`TEST_FRAME_AMOUNT-1) begin
                        PSNR_total = 10*$log10((255.0**2)/($itor(SAD_total)/(3072.0*(`TEST_FRAME_AMOUNT))));
                        
                        if (PSNR_total < `PSNR_BASELINE) begin
                            $display("================ Failed... Your total PSNR = %f, smaller than the required PSNR 23; total latency = %f ns ================\n", PSNR_total, $itor(latency_period_count)*`PERIOD);
                            you_failed_image;
                        end else begin
                            $display("================ Congratulate !!! Your total PSNR = %f, higher that the required PSNR 23; total latency = %f ns ================", PSNR_total, $itor(latency_period_count)*`PERIOD);
                            you_pass_image;
                        end
                        $finish;
                    end
                end

            end
        end
    end


    initial begin
        latency_period_count = 0;

        @(negedge clk);
        while(busy || ~pixel_valid) begin // first input success
            @(negedge clk);
        end

        while(1) begin
            @(negedge clk);
            latency_period_count = latency_period_count + 1;
        end
    end

    initial begin
        repeat(`MAX_LATENCY)@(negedge clk);
        you_failed_image;
        $display("-----------------------------------------------------\n");
        $display("Error!!! The simulation can't be terminated under normal operation!\n");
        $display("-------------------------FAIL------------------------\n");
        $display("-----------------------------------------------------\n");
        $finish;
    end


    always@(negedge clk) begin
        if (ans_frame_count>pat_frame_count) begin
            you_failed_image;
            $display("-----------------------------------------------------\n");
            $display("You cheat !!! You piece of shit !!! It's impossible to output frame %d answer before having %d frame\n", ans_frame_count, pat_frame_count);
            $display("-------------------------FAIL------------------------\n");
            $display("-----------------------------------------------------\n");
            $finish;
        end
    end


    task you_failed_image;
    begin
        $display("\033[38;2;0;0;0m                         \033[38;2;21;22;17m \033[38;2;47;45;41m.\033[38;2;109;106;95m=\033[38;2;119;114;108m=\033[38;2;252;251;247m@\033[38;2;253;254;252m@\033[38;2;252;249;246m@\033[38;2;206;194;183m#\033[38;2;191;173;163m*\033[38;2;176;163;150m*\033[38;2;199;188;169m#\033[38;2;212;196;174m#\033[38;2;107;89;66m-\033[38;2;56;33;2m.\033[38;2;65;46;35m.\033[38;2;19;0;0m \033[38;2;21;6;6m \033[38;2;17;5;1m  \033[38;2;22;1;0m \033[38;2;60;34;21m.\033[38;2;184;173;161m*\033[38;2;201;182;183m#\033[38;2;176;163;162m*\033[38;2;116;97;94m-\033[38;2;87;57;59m:\033[38;2;138;111;101m=\033[38;2;122;103;90m=\033[38;2;83;53;27m:\033[38;2;70;24;1m.\033[38;2;60;6;0m \033[38;2;44;11;1m \033[38;2;76;42;28m.\033[38;2;106;69;50m--\033[38;2;88;47;24m:\033[38;2;57;13;0m \033[38;2;62;30;9m.\033[38;2;29;5;0m \033[38;2;21;16;7m \033[38;2;2;1;4m \033[38;2;1;6;0m \033[38;2;2;10;2m \033[38;2;1;11;3m \033[38;2;0;6;0m  \033[38;2;5;19;3m \033[38;2;9;14;6m \033[38;2;6;16;5m \033[38;2;3;4;4m \033[38;2;1;1;0m \033[38;2;2;2;2m \033[38;2;6;11;4m \033[38;2;24;31;13m.\033[38;2;43;48;26m.\033[38;2;38;41;22m.\033[38;2;57;60;40m:\033[38;2;13;17;4m \033[38;2;11;16;2m \033[38;2;8;11;3m \033[38;2;0;3;2m \033[38;2;10;12;9m \033[38;2;1;1;2m \033[38;2;40;40;33m.\033[38;2;114;117;100m=\033[38;2;205;202;190m#\033[38;2;128;117;115m=\033[38;2;98;79;83m-\033[38;2;58;45;53m.\033[38;2;162;154;159m*\033[38;2;231;226;229m&\033[38;2;139;127;131m+\033[38;2;20;11;14m \033[38;2;8;3;5m \033[38;2;34;25;27m.\033[38;2;71;56;58m:\033[38;2;103;88;89m-\033[38;2;52;37;40m..\033[38;2;14;1;1m \033[38;2;24;2;3m \033[38;2;29;12;5m \033[38;2;53;1;0m \033[38;2;102;36;21m:\033[38;2;127;44;13m:\033[38;2;137;51;4m:\033[38;2;166;94;62m=\033[38;2;152;71;20m-\033[38;2;171;94;71m=\033[38;2;167;90;54m=\033[38;2;204;133;106m+\033[38;2;193;130;112m+\033[38;2;220;154;131m*\033[38;2;221;166;143m*\033[0m");
        $display("\033[38;2;0;0;0m                       \033[38;2;33;30;42m.\033[38;2;48;42;57m.\033[38;2;214;210;210m&\033[38;2;254;253;253m@\033[38;2;245;236;239m@\033[38;2;254;254;252m@\033[38;2;248;241;238m@\033[38;2;255;249;242m@\033[38;2;226;204;201m&\033[38;2;240;221;223m&\033[38;2;249;239;239m@\033[38;2;255;251;254m@@\033[38;2;141;128;120m+\033[38;2;158;139;129m+\033[38;2;121;101;76m=\033[38;2;52;24;17m.\033[38;2;125;107;91m=\033[38;2;31;19;6m \033[38;2;18;11;4m  \033[38;2;31;7;2m \033[38;2;37;4;0m \033[38;2;149;133;123m+\033[38;2;229;215;215m&\033[38;2;175;154;155m*\033[38;2;132;98;98m=\033[38;2;58;21;20m.\033[38;2;56;31;8m.\033[38;2;33;1;0m   \033[38;2;93;44;26m:\033[38;2;99;62;40m:\033[38;2;117;96;77m-\033[38;2;114;81;66m-\033[38;2;48;22;5m.\033[38;2;91;57;49m:\033[38;2;168;134;113m+\033[38;2;192;169;149m*\033[38;2;112;88;42m-\033[38;2;114;91;59m-\033[38;2;54;37;20m.\033[38;2;24;22;10m \033[38;2;12;18;8m \033[38;2;4;13;2m \033[38;2;3;17;4m \033[38;2;2;20;1m \033[38;2;39;59;30m.\033[38;2;228;229;215m&\033[38;2;146;154;131m+\033[38;2;19;21;10m \033[38;2;10;13;1m  \033[38;2;5;11;4m \033[38;2;4;18;3m \033[38;2;3;15;1m \033[38;2;1;11;2m \033[38;2;7;9;5m \033[38;2;1;4;1m   \033[38;2;10;13;6m \033[38;2;3;10;0m \033[38;2;32;29;16m.\033[38;2;95;84;78m-\033[38;2;133;127;116m=\033[38;2;80;70;59m:\033[38;2;26;9;5m \033[38;2;40;18;19m  \033[38;2;193;186;181m#\033[38;2;172;156;155m*\033[38;2;22;18;14m \033[38;2;20;10;8m \033[38;2;14;1;1m \033[38;2;54;37;34m.\033[38;2;53;30;27m.\033[38;2;36;17;14m \033[38;2;42;24;24m.\033[38;2;20;0;1m \033[38;2;24;6;2m  \033[38;2;56;15;13m.\033[38;2;100;37;36m:\033[38;2;127;62;33m-\033[38;2;151;84;50m-\033[38;2;149;73;34m-\033[38;2;136;56;10m:\033[38;2;172;90;53m=\033[38;2;165;93;59m=\033[38;2;209;137;109m+\033[38;2;196;131;104m+\033[38;2;214;157;130m*\033[38;2;203;140;115m*\033[38;2;216;163;138m*\033[0m");
        $display("\033[38;2;0;0;0m                    \033[38;2;2;2;4m \033[38;2;13;12;18m \033[38;2;59;56;67m:\033[38;2;171;167;182m*\033[38;2;255;254;253m@@@@\033[38;2;178;155;142m*\033[38;2;242;219;206m&\033[38;2;195;178;164m*\033[38;2;253;252;238m@\033[38;2;247;235;232m@\033[38;2;254;250;249m@\033[38;2;255;253;251m@\033[38;2;245;234;229m@\033[38;2;206;182;178m#\033[38;2;252;252;248m@\033[38;2;230;210;203m&\033[38;2;243;236;229m@\033[38;2;74;55;41m:\033[38;2;38;15;7m \033[38;2;29;1;6m  \033[38;2;115;76;63m-\033[38;2;63;14;6m.\033[38;2;61;5;0m \033[38;2;101;52;34m:\033[38;2;111;51;43m:\033[38;2;101;46;34m:\033[38;2;84;22;7m.\033[38;2;117;72;45m-\033[38;2;74;29;1m.\033[38;2;89;22;13m.\033[38;2;59;1;0m \033[38;2;55;0;6m \033[38;2;35;3;0m \033[38;2;59;39;11m.\033[38;2;57;27;4m.\033[38;2;61;24;18m.\033[38;2;106;54;55m:\033[38;2;69;23;20m.\033[38;2;54;1;1m \033[38;2;125;88;59m-\033[38;2;161;139;111m+\033[38;2;112;88;47m-\033[38;2;107;80;50m-\033[38;2;35;23;3m \033[38;2;30;19;8m \033[38;2;6;0;0m \033[38;2;2;7;1m \033[38;2;6;12;0m \033[38;2;101;106;87m-\033[38;2;22;26;9m \033[38;2;12;16;1m \033[38;2;7;7;4m \033[38;2;3;4;3m \033[38;2;1;0;0m \033[38;2;4;11;3m \033[38;2;3;16;5m \033[38;2;2;14;2m  \033[38;2;0;7;1m \033[38;2;3;25;6m \033[38;2;0;17;1m \033[38;2;3;9;0m  \033[38;2;105;99;85m-\033[38;2;224;215;208m&\033[38;2;23;9;1m \033[38;2;22;4;2m \033[38;2;32;15;13m \033[38;2;15;2;0m \033[38;2;86;73;65m:\033[38;2;108;91;87m-\033[38;2;23;2;3m \033[38;2;13;0;2m \033[38;2;17;1;1m \033[38;2;18;3;4m \033[38;2;25;7;7m \033[38;2;22;0;2m \033[38;2;16;2;1m \033[38;2;24;1;3m  \033[38;2;22;4;2m \033[38;2;35;0;0m  \033[38;2;136;70;54m-\033[38;2;131;63;28m-\033[38;2;120;32;0m:\033[38;2;150;70;28m--\033[38;2;175;99;62m==\033[38;2;171;93;45m=\033[38;2;163;87;46m=\033[38;2;185;116;85m+\033[38;2;172;105;62m=\033[38;2;185;127;96m+\033[0m");
        $display("\033[38;2;0;0;0m                 \033[38;2;5;5;5m \033[38;2;1;1;1m  \033[38;2;30;27;28m.\033[38;2;96;95;100m-\033[38;2;253;251;253m@\033[38;2;252;250;254m@@\033[38;2;255;252;245m@\033[38;2;247;237;227m@\033[38;2;168;143;118m+\033[38;2;232;203;187m&\033[38;2;122;97;54m-\033[38;2;206;192;168m#\033[38;2;209;189;172m#\033[38;2;239;237;222m@\033[38;2;243;231;216m&\033[38;2;154;132;111m+\033[38;2;100;58;28m:\033[38;2;189;156;132m*\033[38;2;148;124;77m=\033[38;2;103;81;13m-\033[38;2;61;25;3m.\033[38;2;60;1;6m \033[38;2;85;24;11m.\033[38;2;76;21;2m.\033[38;2;111;49;31m:\033[38;2;140;86;59m-\033[38;2;115;54;27m:\033[38;2;150;104;79m=\033[38;2;180;131;114m+\033[38;2;164;107;74m=\033[38;2;178;116;102m+\033[38;2;154;90;74m=\033[38;2;170;104;83m=\033[38;2;190;125;109m+\033[38;2;178;120;104m+\033[38;2;171;124;98m+\033[38;2;168;113;97m=\033[38;2;160;114;87m=\033[38;2;164;116;99m=\033[38;2;178;131;107m+\033[38;2;124;61;52m-\033[38;2;67;3;0m \033[38;2;55;1;3m  \033[38;2;93;28;28m.\033[38;2;50;1;1m \033[38;2;194;163;132m*\033[38;2;141;112;85m=\033[38;2;119;79;58m-\033[38;2;82;40;16m.\033[38;2;66;45;38m.\033[38;2;4;1;4m \033[38;2;2;0;3m \033[38;2;0;7;0m \033[38;2;10;16;2m \033[38;2;5;8;1m \033[38;2;4;1;2m  \033[38;2;5;7;4m  \033[38;2;0;2;0m \033[38;2;4;14;7m  \033[38;2;1;1;1m   \033[38;2;7;15;0m \033[38;2;28;26;13m \033[38;2;75;71;58m:\033[38;2;17;3;0m \033[38;2;22;5;1m  \033[38;2;14;6;4m \033[38;2;38;25;20m.\033[38;2;32;15;8m \033[38;2;67;57;55m:\033[38;2;20;5;5m \033[38;2;12;1;1m  \033[38;2;20;3;4m \033[38;2;13;1;0m  \033[38;2;22;2;3m  \033[38;2;21;7;6m \033[38;2;26;0;1m  \033[38;2;120;70;62m-\033[38;2;141;83;64m-\033[38;2;126;60;35m:\033[38;2;130;66;22m-\033[38;2;158;92;59m=\033[38;2;160;96;62m=\033[38;2;152;82;44m-\033[38;2;164;90;59m=\033[38;2;160;80;33m-\033[38;2;179;110;74m=\033[38;2;195;131;102m+\033[38;2;186;121;93m+\033[38;2;211;157;133m*\033[0m");
        $display("\033[38;2;0;0;0m                 \033[38;2;7;4;5m \033[38;2;26;19;12m \033[38;2;94;89;98m-\033[38;2;243;238;244m@\033[38;2;253;253;255m@\033[38;2;255;254;252m@\033[38;2;240;232;227m@\033[38;2;255;253;244m@\033[38;2;248;228;214m&\033[38;2;159;131;87m+\033[38;2;210;179;151m#\033[38;2;126;79;47m-\033[38;2;167;133;102m+\033[38;2;210;182;155m#\033[38;2;218;195;170m#\033[38;2;249;236;212m@\033[38;2;183;160;126m*\033[38;2;150;115;72m=\033[38;2;105;54;5m:\033[38;2;192;156;132m*\033[38;2;133;92;39m-\033[38;2;157;97;62m=\033[38;2;117;47;2m:\033[38;2;172;119;80m+\033[38;2;130;64;13m-\033[38;2;158;98;63m=\033[38;2;178;123;89m+\033[38;2;186;121;94m+\033[38;2;184;120;93m+\033[38;2;183;114;84m+\033[38;2;182;112;80m=\033[38;2;185;124;98m+\033[38;2;184;114;83m++\033[38;2;193;123;100m+\033[38;2;188;122;96m+\033[38;2;189;121;100m+\033[38;2;194;123;103m+\033[38;2;183;108;80m=\033[38;2;178;107;84m=\033[38;2;171;100;78m=\033[38;2;177;104;83m=\033[38;2;163;89;72m=\033[38;2;165;99;82m=\033[38;2;162;113;90m=\033[38;2;130;63;56m-\033[38;2;71;3;1m \033[38;2;61;0;2m \033[38;2;86;18;17m.\033[38;2;101;45;33m:\033[38;2;173;138;111m+\033[38;2;130;94;69m-\033[38;2;71;44;6m.\033[38;2;32;12;1m  \033[38;2;10;9;5m \033[38;2;3;0;0m    \033[38;2;1;1;1m  \033[38;2;2;16;3m \033[38;2;3;13;2m \033[38;2;9;18;6m \033[38;2;5;14;4m \033[38;2;0;3;1m \033[38;2;1;1;3m \033[38;2;5;5;0m \033[38;2;44;39;33m.\033[38;2;29;9;6m \033[38;2;26;0;0m    \033[38;2;44;27;19m..\033[38;2;21;2;1m  \033[38;2;9;1;0m \033[38;2;38;2;4m \033[38;2;11;0;0m    \033[38;2;20;4;4m \033[38;2;26;0;3m  \033[38;2;35;3;0m \033[38;2;45;10;2m  \033[38;2;53;25;4m.\033[38;2;55;28;7m.\033[38;2;69;39;21m.\033[38;2;50;21;6m.\033[38;2;65;41;25m.\033[38;2;47;8;8m \033[38;2;52;1;1m \033[38;2;116;31;22m:\033[38;2;202;145;114m*\033[38;2;198;138;108m+\033[38;2;202;145;125m*\033[0m");
        $display("\033[38;2;0;0;0m                 \033[38;2;7;5;4m \033[38;2;52;44;38m.\033[38;2;254;251;251m@\033[38;2;253;254;249m@\033[38;2;211;192;181m#\033[38;2;234;213;200m&&\033[38;2;244;229;210m&\033[38;2;158;129;85m+\033[38;2;176;154;113m*\033[38;2;166;136;101m+\033[38;2;119;66;28m-\033[38;2;252;230;218m@\033[38;2;208;189;167m#\033[38;2;250;234;208m@\033[38;2;134;76;51m-\033[38;2;195;169;143m*\033[38;2;106;51;40m:\033[38;2;143;93;61m=\033[38;2;206;175;147m*\033[38;2;134;74;20m-\033[38;2;177;109;88m=\033[38;2;172;113;85m=\033[38;2;139;64;13m-\033[38;2;173;103;75m=\033[38;2;180;119;83m+\033[38;2;196;125;99m+\033[38;2;199;124;105m+\033[38;2;189;118;95m+\033[38;2;210;144;120m*\033[38;2;189;123;100m+\033[38;2;174;98;62m=\033[38;2;194;122;99m+\033[38;2;186;120;89m+\033[38;2;192;124;102m+\033[38;2;203;135;112m++\033[38;2;199;131;110m+\033[38;2;195;127;106m+\033[38;2;190;123;97m+\033[38;2;177;103;75m=\033[38;2;182;106;82m==\033[38;2;166;92;67m=\033[38;2;175;105;84m=\033[38;2;172;95;69m=\033[38;2;200;142;126m*\033[38;2;183;124;106m+\033[38;2;98;6;10m.\033[38;2;60;1;3m \033[38;2;89;10;9m.\033[38;2;217;179;167m#\033[38;2;172;140;114m+\033[38;2;121;90;67m-\033[38;2;36;2;0m   \033[38;2;0;0;2m   \033[38;2;1;1;1m \033[38;2;2;4;0m \033[38;2;1;16;3m \033[38;2;4;15;0m \033[38;2;14;24;12m \033[38;2;4;8;2m \033[38;2;2;1;4m \033[38;2;1;3;2m \033[38;2;15;8;6m \033[38;2;20;4;5m  \033[38;2;15;0;4m   \033[38;2;18;3;0m \033[38;2;14;7;1m \033[38;2;20;1;3m \033[38;2;8;0;0m   \033[38;2;19;2;2m  \033[38;2;26;0;0m   \033[38;2;29;2;5m \033[38;2;28;0;3m \033[38;2;47;22;20m.\033[38;2;100;67;61m:\033[38;2;101;63;53m:\033[38;2;102;59;48m:\033[38;2;125;86;71m-\033[38;2;158;134;120m+\033[38;2;97;69;60m:\033[38;2;75;45;39m:\033[38;2;35;6;0m  \033[38;2;47;13;3m \033[38;2;62;2;1m \033[38;2;89;0;3m.\033[38;2;168;98;75m=\033[38;2;180;118;92m+\033[0m");
        $display("\033[38;2;0;0;0m                \033[38;2;7;7;7m \033[38;2;31;27;23m.\033[38;2;252;247;242m@\033[38;2;249;252;248m@\033[38;2;205;178;171m#\033[38;2;201;170;144m*\033[38;2;228;205;176m&\033[38;2;229;214;198m&\033[38;2;140;116;87m=\033[38;2;104;44;32m:\033[38;2;231;215;195m&\033[38;2;128;79;71m-\033[38;2;217;187;169m#\033[38;2;207;180;157m#\033[38;2;251;236;225m@\033[38;2;243;206;191m&\033[38;2;143;89;58m-\033[38;2;156;124;81m=\033[38;2;100;39;24m:\033[38;2;149;97;65m=\033[38;2;183;142;124m+\033[38;2;126;58;31m:\033[38;2;174;118;94m+\033[38;2;170;95;72m=\033[38;2;187;111;87m+\033[38;2;193;123;97m++\033[38;2;202;119;98m++\033[38;2;188;106;82m=\033[38;2;206;136;111m+\033[38;2;187;111;79m+\033[38;2;216;149;129m**\033[38;2;195;126;97m+\033[38;2;192;123;94m+\033[38;2;197;126;105m+\033[38;2;194;127;101m+\033[38;2;198;131;105m+\033[38;2;211;148;124m*\033[38;2;212;146;120m*\033[38;2;182;107;78m=\033[38;2;173;100;70m=\033[38;2;191;125;99m+\033[38;2;204;143;122m*\033[38;2;188;117;92m+\033[38;2;160;70;42m-\033[38;2;172;93;61m=\033[38;2;167;103;80m=\033[38;2;170;110;79m=\033[38;2;145;62;48m-\033[38;2;87;0;1m.\033[38;2;103;22;2m.\033[38;2;197;162;129m*\033[38;2;218;188;160m#\033[38;2;127;85;62m-\033[38;2;41;23;5m. \033[38;2;1;1;3m \033[38;2;0;0;0m  \033[38;2;1;1;1m    \033[38;2;0;9;2m \033[38;2;6;15;4m \033[38;2;29;27;22m.\033[38;2;19;20;14m \033[38;2;16;2;1m \033[38;2;22;1;2m \033[38;2;25;0;3m  \033[38;2;26;2;2m \033[38;2;20;1;0m  \033[38;2;29;0;4m    \033[38;2;26;1;1m  \033[38;2;28;2;3m \033[38;2;12;0;0m  \033[38;2;31;1;1m  \033[38;2;19;0;0m  \033[38;2;31;1;1m \033[38;2;34;4;0m \033[38;2;76;50;41m:\033[38;2;125;98;87m=\033[38;2;170;145;135m+\033[38;2;173;141;134m+\033[38;2;126;87;81m-\033[38;2;63;19;20m.\033[38;2;44;1;1m \033[38;2;74;19;4m.\033[38;2;110;43;27m:\033[38;2;140;77;47m-\033[38;2;161;97;62m=\033[38;2;187;137;111m+\033[0m");
        $display("\033[38;2;0;0;0m             \033[38;2;1;1;1m   \033[38;2;59;57;44m:\033[38;2;243;233;224m@\033[38;2;252;246;245m@\033[38;2;250;229;203m&\033[38;2;217;183;155m#\033[38;2;225;200;177m#\033[38;2;242;219;202m&\033[38;2;230;218;205m&\033[38;2;74;4;2m \033[38;2;186;142;121m+\033[38;2;247;218;203m&\033[38;2;162;117;86m=\033[38;2;217;185;159m#\033[38;2;194;153;112m*\033[38;2;252;252;244m@\033[38;2;123;72;47m-\033[38;2;206;177;153m#\033[38;2;127;84;16m-\033[38;2;124;61;2m:\033[38;2;173;132;96m+\033[38;2;153;85;64m-\033[38;2;169;104;77m=\033[38;2;154;92;39m=\033[38;2;161;81;16m-\033[38;2;198;124;95m+\033[38;2;180;109;84m=\033[38;2;195;120;95m+\033[38;2;203;126;105m+\033[38;2;221;150;132m*\033[38;2;214;146;127m*\033[38;2;210;139;119m*\033[38;2;211;142;122m*\033[38;2;210;139;119m*\033[38;2;206;135;115m+\033[38;2;203;132;112m+\033[38;2;211;140;120m*\033[38;2;217;146;126m*\033[38;2;209;138;118m*\033[38;2;210;139;119m*\033[38;2;219;148;130m*\033[38;2;211;143;124m*\033[38;2;200;133;114m+\033[38;2;212;144;125m*\033[38;2;187;115;97m+\033[38;2;201;132;116m+\033[38;2;187;119;100m+\033[38;2;173;103;77m=\033[38;2;185;114;92m+\033[38;2;197;130;112m+\033[38;2;183;110;93m+\033[38;2;165;94;64m=\033[38;2;188;116;95m+\033[38;2;101;23;9m.\033[38;2;77;0;1m \033[38;2;141;73;38m-\033[38;2;237;208;183m&\033[38;2;127;99;65m-\033[38;2;80;54;32m:\033[38;2;20;10;11m \033[38;2;2;1;2m  \033[38;2;0;0;0m   \033[38;2;1;1;1m \033[38;2;7;9;5m \033[38;2;78;82;75m-\033[38;2;9;9;4m \033[38;2;6;1;0m \033[38;2;14;4;3m  \033[38;2;3;1;2m   \033[38;2;0;0;0m     \033[38;2;1;1;1m \033[38;2;0;2;4m  \033[38;2;6;0;2m \033[38;2;29;2;5m \033[38;2;37;0;4m \033[38;2;20;1;2m \033[38;2;39;20;17m \033[38;2;28;2;3m \033[38;2;3;0;1m  \033[38;2;29;4;3m \033[38;2;48;24;20m.\033[38;2;90;69;62m:\033[38;2;66;47;40m:\033[38;2;23;6;4m \033[38;2;35;1;7m \033[38;2;45;5;5m \033[38;2;40;1;0m \033[38;2;65;9;12m.\033[38;2;67;1;2m \033[38;2;95;19;5m.\033[38;2;108;20;1m.\033[38;2;174;117;91m+\033[0m");
        $display("\033[38;2;0;0;0m              \033[38;2;9;17;14m \033[38;2;46;38;22m.\033[38;2;215;207;182m#\033[38;2;212;195;179m#\033[38;2;253;239;221m@\033[38;2;254;228;202m&\033[38;2;226;201;170m#\033[38;2;197;167;137m*\033[38;2;246;233;211m@\033[38;2;61;6;0m \033[38;2;165;130;100m+\033[38;2;201;173;147m*\033[38;2;188;160;129m*\033[38;2;226;194;167m#\033[38;2;124;72;16m-\033[38;2;212;183;153m#\033[38;2;252;248;238m@\033[38;2;85;10;5m.\033[38;2;199;167;147m*\033[38;2;191;149;100m*\033[38;2;133;63;11m-\033[38;2;196;153;111m*\033[38;2;141;71;25m-\033[38;2;203;139;105m+\033[38;2;172;107;66m==\033[38;2;226;156;131m*\033[38;2;215;144;123m*\033[38;2;217;141;116m*\033[38;2;194;113;86m+\033[38;2;213;142;122m*\033[38;2;227;159;138m*\033[38;2;215;142;123m*\033[38;2;211;140;120m*\033[38;2;206;135;115m+\033[38;2;218;150;129m***\033[38;2;228;157;137m*\033[38;2;226;159;140m**\033[38;2;229;162;143m*\033[38;2;225;156;140m*\033[38;2;236;171;153m#\033[38;2;207;141;124m*\033[38;2;211;142;126m*\033[38;2;224;160;143m*\033[38;2;237;174;157m#\033[38;2;214;147;128m*\033[38;2;178;110;89m=\033[38;2;193;125;106m+\033[38;2;183;112;92m+\033[38;2;182;106;86m=\033[38;2;176;107;84m=\033[38;2;173;108;87m=\033[38;2;163;93;68m=\033[38;2;69;1;0m \033[38;2;164;107;82m=\033[38;2;176;149;112m+\033[38;2;145;115;87m=\033[38;2;58;37;17m.\033[38;2;4;3;4m  \033[38;2;2;0;1m   \033[38;2;1;12;4m \033[38;2;3;17;6m \033[38;2;1;6;1m \033[38;2;7;8;4m \033[38;2;21;14;11m \033[38;2;7;3;4m \033[38;2;1;1;1m \033[38;2;0;0;0m     \033[38;2;1;1;1m      \033[38;2;35;2;5m \033[38;2;36;0;0m \033[38;2;31;10;5m \033[38;2;28;11;4m \033[38;2;31;5;2m \033[38;2;37;4;0m \033[38;2;44;9;5m \033[38;2;29;7;0m \033[38;2;55;16;10m.\033[38;2;83;50;40m:\033[38;2;138;104;94m=\033[38;2;44;16;11m \033[38;2;32;7;2m \033[38;2;43;10;6m \033[38;2;83;56;53m:\033[38;2;39;1;0m \033[38;2;78;32;26m.\033[38;2;67;2;2m \033[38;2;79;0;1m \033[38;2;86;6;0m.\033[38;2;159;105;74m=\033[0m");
        $display("\033[38;2;0;0;0m             \033[38;2;17;17;9m \033[38;2;29;12;0m \033[38;2;172;152;132m*\033[38;2;159;137;106m+\033[38;2;251;242;228m@\033[38;2;240;216;194m&\033[38;2;238;214;182m&\033[38;2;209;177;145m#\033[38;2;231;209;185m&\033[38;2;174;134;110m+\033[38;2;125;66;24m-\033[38;2;190;168;121m*\033[38;2;255;236;203m@\033[38;2;192;164;132m*\033[38;2;186;149;97m+\033[38;2;146;96;44m=\033[38;2;254;242;218m@\033[38;2;250;239;216m@\033[38;2;75;5;3m.\033[38;2;197;168;139m*\033[38;2;234;201;170m#\033[38;2;145;80;5m-\033[38;2;206;165;121m**\033[38;2;227;176;148m#\033[38;2;165;93;37m=\033[38;2;164;74;20m-\033[38;2;213;141;109m*\033[38;2;186;116;87m+\033[38;2;212;135;105m+\033[38;2;196;121;82m+\033[38;2;216;139;109m*\033[38;2;221;149;124m*\033[38;2;224;156;136m*\033[38;2;219;151;132m*\033[38;2;243;178;160m#\033[38;2;240;173;157m#\033[38;2;246;178;164m#\033[38;2;223;158;140m*\033[38;2;225;164;146m*\033[38;2;238;176;161m##\033[38;2;228;168;150m#\033[38;2;217;152;134m*\033[38;2;209;144;124m*\033[38;2;220;154;136m*\033[38;2;213;149;131m*\033[38;2;200;132;113m+\033[38;2;204;139;121m*\033[38;2;228;162;146m*\033[38;2;200;133;115m+\033[38;2;192;121;93m+\033[38;2;209;144;124m*\033[38;2;187;111;96m+\033[38;2;173;101;74m=\033[38;2;165;94;62m=\033[38;2;181;121;93m+\033[38;2;103;18;6m.\033[38;2;86;7;3m.\033[38;2;143;91;62m-\033[38;2;159;119;86m=\033[38;2;134;107;81m=\033[38;2;35;20;5m \033[38;2;2;0;3m \033[38;2;0;1;0m        \033[38;2;2;0;1m             \033[38;2;38;2;4m \033[38;2;35;3;1m \033[38;2;43;2;3m \033[38;2;67;3;1m \033[38;2;113;64;48m:\033[38;2;128;73;52m-\033[38;2;101;45;9m:\033[38;2;135;86;73m-\033[38;2;130;78;69m-\033[38;2;83;18;10m.\033[38;2;77;2;6m \033[38;2;85;18;1m.\033[38;2;100;37;11m:\033[38;2;97;24;10m.\033[38;2;90;14;2m.\033[38;2;108;48;30m:\033[38;2;94;25;10m.\033[38;2;71;2;2m \033[38;2;62;1;0m \033[38;2;98;20;7m.\033[38;2;129;66;38m-\033[0m");
        $display("\033[38;2;0;0;0m             \033[38;2;60;55;37m:\033[38;2;119;92;67m-\033[38;2;211;187;165m#\033[38;2;192;163;128m*\033[38;2;251;227;213m&\033[38;2;245;215;185m&\033[38;2;224;195;157m#\033[38;2;197;166;133m*\033[38;2;248;228;206m&\033[38;2;102;39;24m:\033[38;2;177;134;96m+\033[38;2;218;188;163m#\033[38;2;229;211;179m&\033[38;2;237;209;174m&\033[38;2;154;113;51m=\033[38;2;223;182;147m#\033[38;2;254;232;202m@\033[38;2;255;246;227m@\033[38;2;78;8;1m.\033[38;2;127;59;43m-\033[38;2;241;221;200m&\033[38;2;137;56;1m:\033[38;2;209;166;123m*\033[38;2;182;121;70m+\033[38;2;233;192;156m#\033[38;2;189;115;78m+\033[38;2;212;149;114m*\033[38;2;222;154;125m*\033[38;2;207;138;107m+\033[38;2;220;149;123m*\033[38;2;200;130;98m+\033[38;2;209;138;113m*\033[38;2;230;162;141m*\033[38;2;236;170;153m#\033[38;2;250;185;166m#\033[38;2;230;165;147m#\033[38;2;234;172;152m#\033[38;2;239;175;158m#\033[38;2;232;166;148m#\033[38;2;224;159;140m*\033[38;2;202;134;115m+\033[38;2;206;135;120m+\033[38;2;208;137;127m*\033[38;2;237;183;167m#\033[38;2;238;180;164m#\033[38;2;200;138;120m+\033[38;2;210;142;122m*\033[38;2;201;132;112m+\033[38;2;206;133;115m+\033[38;2;192;125;103m+\033[38;2;211;146;123m*\033[38;2;175;98;75m=\033[38;2;160;88;63m=\033[38;2;190;122;97m+\033[38;2;180;114;85m+\033[38;2;165;100;73m=\033[38;2;203;137;110m+\033[38;2;189;135;106m+\033[38;2;104;35;19m:\033[38;2;63;1;4m \033[38;2;110;66;30m:\033[38;2;139;106;75m=\033[38;2;162;142;112m+\033[38;2;62;52;35m:\033[38;2;1;1;0m \033[38;2;0;0;1m                  \033[38;2;3;1;2m \033[38;2;21;3;5m \033[38;2;37;0;2m \033[38;2;48;15;9m \033[38;2;92;22;20m.\033[38;2;126;72;47m-\033[38;2;151;95;67m=\033[38;2;134;62;32m-\033[38;2;125;59;18m:\033[38;2;160;100;67m=\033[38;2;182;124;104m+\033[38;2;147;87;58m-\033[38;2;145;82;49m-\033[38;2;148;84;43m-\033[38;2;160;100;72m=\033[38;2;163;105;80m=\033[38;2;153;95;74m=\033[38;2;148;91;81m=\033[38;2;112;46;26m:\033[38;2;71;5;3m \033[38;2;87;2;0m.\033[38;2;122;53;32m:\033[38;2;136;74;56m-\033[0m");
        $display("\033[38;2;0;0;0m            \033[38;2;29;33;17m.\033[38;2;53;55;29m.\033[38;2;221;208;188m&\033[38;2;143;100;61m=\033[38;2;245;227;197m&\033[38;2;247;217;190m&\033[38;2;228;190;158m#\033[38;2;215;176;146m#\033[38;2;250;226;203m&\033[38;2;130;74;39m-\033[38;2;121;65;6m:\033[38;2;149;101;37m=\033[38;2;253;238;213m@\033[38;2;142;97;41m=\033[38;2;235;204;170m&\033[38;2;157;104;43m=\033[38;2;233;198;165m#\033[38;2;255;238;212m@\033[38;2;226;187;163m#\033[38;2;95;27;12m.\033[38;2;131;62;55m-\033[38;2;242;227;202m&\033[38;2;165;98;41m=\033[38;2;189;133;81m+\033[38;2;248;220;190m&\033[38;2;210;158;117m*\033[38;2;186;113;62m=\033[38;2;224;159;132m*\033[38;2;225;155;130m*\033[38;2;227;160;132m*\033[38;2;232;164;141m#\033[38;2;227;160;136m*\033[38;2;241;174;153m#\033[38;2;232;165;143m#\033[38;2;224;157;140m*\033[38;2;210;143;124m*\033[38;2;217;144;125m*\033[38;2;213;140;121m**\033[38;2;211;143;124m*\033[38;2;203;135;116m+\033[38;2;197;126;106m+\033[38;2;215;142;125m*\033[38;2;212;144;127m*\033[38;2;188;121;101m+\033[38;2;218;157;139m*\033[38;2;241;181;163m#\033[38;2;220;153;134m****\033[38;2;221;156;139m*\033[38;2;239;190;171m#\033[38;2;184;113;95m+\033[38;2;195;125;104m+\033[38;2;181;133;110m+\033[38;2;208;154;137m*\033[38;2;186;143;119m+\033[38;2;192;140;127m+\033[38;2;175;129;102m+\033[38;2;70;7;8m.\033[38;2;64;5;5m \033[38;2;106;68;42m:\033[38;2;119;72;45m-\033[38;2;157;129;119m+\033[38;2;18;12;4m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m  \033[38;2;7;1;2m  \033[38;2;2;0;1m            \033[38;2;1;1;0m \033[38;2;32;2;4m  \033[38;2;66;4;1m \033[38;2;135;73;55m-\033[38;2;136;65;37m-\033[38;2;150;74;43m-\033[38;2;142;66;24m-\033[38;2;150;77;45m-\033[38;2;147;74;28m-\033[38;2;165;96;60m=\033[38;2;169;107;63m=\033[38;2;178;116;85m+\033[38;2;187;138;102m+\033[38;2;185;134;99m+\033[38;2;198;149;122m*\033[38;2;169;110;85m=\033[38;2;107;29;7m.\033[38;2;76;3;1m \033[38;2;69;0;0m \033[38;2;131;64;45m-\033[38;2;137;73;46m-\033[38;2;139;69;44m-\033[0m");
        $display("\033[38;2;0;0;0m         \033[38;2;1;1;1m  \033[38;2;10;5;2m \033[38;2;48;29;26m.\033[38;2;190;171;165m*\033[38;2;203;163;146m*\033[38;2;191;151;115m*\033[38;2;245;229;209m&\033[38;2;241;214;190m&\033[38;2;209;179;155m#\033[38;2;242;215;185m&\033[38;2;178;131;94m+\033[38;2;72;9;0m.\033[38;2;216;179;156m#\033[38;2;123;52;45m:\033[38;2;217;190;152m#\033[38;2;211;173;119m*\033[38;2;238;191;154m#\033[38;2;141;95;10m-\033[38;2;249;219;197m&\033[38;2;250;222;195m&\033[38;2;209;169;143m*\033[38;2;84;7;8m.\033[38;2;125;48;43m:\033[38;2;255;233;218m@\033[38;2;153;77;4m-\033[38;2;186;130;82m+\033[38;2;255;238;212m@\033[38;2;182;106;48m=\033[38;2;206;137;102m+\033[38;2;218;150;126m*\033[38;2;222;153;124m**\033[38;2;226;158;130m*\033[38;2;228;161;134m*\033[38;2;237;169;148m#\033[38;2;233;165;146m#\033[38;2;231;159;145m**\033[38;2;220;145;129m*\033[38;2;221;147;128m*\033[38;2;215;144;126m*\033[38;2;217;149;132m*\033[38;2;219;156;139m*\033[38;2;231;170;155m#\033[38;2;228;159;144m*\033[38;2;229;155;143m*\033[38;2;211;144;127m*\033[38;2;207;137;121m*\033[38;2;223;157;142m*\033[38;2;245;187;171m#\033[38;2;250;188;173m#\033[38;2;238;178;169m#\033[38;2;222;162;143m*\033[38;2;233;173;159m#\033[38;2;253;225;207m&\033[38;2;209;155;134m*\033[38;2;106;40;24m:\033[38;2;63;2;1m \033[38;2;47;0;2m \033[38;2;53;4;10m \033[38;2;52;1;2m \033[38;2;53;2;0m \033[38;2;78;24;21m.\033[38;2;42;1;2m \033[38;2;78;5;4m.\033[38;2;105;49;24m:\033[38;2;134;103;74m=\033[38;2;125;104;78m=\033[38;2;42;23;9m.\033[38;2;3;1;5m   \033[38;2;16;11;9m \033[38;2;12;2;2m  \033[38;2;2;0;1m           \033[38;2;38;1;0m  \033[38;2;75;26;5m.\033[38;2;92;17;0m.\033[38;2;93;3;2m.\033[38;2;118;34;0m:\033[38;2;133;52;6m:\033[38;2;139;60;7m-:\033[38;2;156;71;28m-\033[38;2;172;99;65m=\033[38;2;184;111;85m+\033[38;2;178;112;81m=\033[38;2;181;105;75m=\033[38;2;174;98;71m=\033[38;2;181;117;89m+\033[38;2;139;62;37m-\033[38;2;74;3;2m \033[38;2;66;4;4m \033[38;2;196;141;142m*+\033[38;2;120;37;12m:\033[38;2;135;65;47m-\033[0m");
        $display("\033[38;2;0;0;0m           \033[38;2;37;31;20m.\033[38;2;106;88;75m-\033[38;2;197;173;157m*\033[38;2;101;44;4m:\033[38;2;250;227;205m&\033[38;2;249;225;195m&\033[38;2;232;200;175m#\033[38;2;213;182;155m#\033[38;2;190;153;122m*\033[38;2;142;106;49m=\033[38;2;157;117;82m=\033[38;2;88;24;15m.\033[38;2;249;219;183m&\033[38;2;156;107;48m=\033[38;2;232;198;161m#\033[38;2;142;94;18m-\033[38;2;199;156;117m*\033[38;2;255;230;209m@\033[38;2;188;138;105m+\033[38;2;237;194;172m#\033[38;2;82;0;3m \033[38;2;154;81;58m-\033[38;2;252;233;215m@\033[38;2;139;58;3m:\033[38;2;219;174;128m#\033[38;2;252;239;220m@\033[38;2;149;71;32m-\033[38;2;220;150;125m**\033[38;2;230;166;138m#\033[38;2;227;163;135m*\033[38;2;222;162;133m*\033[38;2;236;176;149m#\033[38;2;240;180;156m#\033[38;2;233;167;151m#\033[38;2;239;172;152m#\033[38;2;220;156;134m*\033[38;2;235;178;153m#\033[38;2;242;191;174m#\033[38;2;254;214;201m&\033[38;2;245;198;183m&\033[38;2;255;210;192m&\033[38;2;239;184;170m#\033[38;2;255;204;190m&&\033[38;2;248;195;181m&\033[38;2;232;166;151m#\033[38;2;218;157;138m*\033[38;2;240;178;165m##\033[38;2;206;136;123m+\033[38;2;222;156;139m*\033[38;2;155;84;58m-\033[38;2;78;4;1m.\033[38;2;47;0;4m    \033[38;2;117;62;45m:\033[38;2;173;123;98m+\033[38;2;182;138;120m+\033[38;2;217;185;163m#\033[38;2;122;74;65m-\033[38;2;89;45;42m:\033[38;2;60;0;0m \033[38;2;117;64;34m:\033[38;2;153;119;92m=\033[38;2;115;89;67m-\033[38;2;38;30;16m.\033[38;2;20;13;3m \033[38;2;9;4;1m \033[38;2;23;7;8m \033[38;2;6;1;1m  \033[38;2;9;0;3m \033[38;2;1;1;1m \033[38;2;0;0;0m          \033[38;2;56;12;9m \033[38;2;72;11;8m.\033[38;2;94;13;4m.\033[38;2;100;18;10m.\033[38;2;110;8;4m.\033[38;2;104;5;0m.\033[38;2;129;39;4m:\033[38;2;152;69;34m-\033[38;2;170;98;72m=\033[38;2;161;87;49m=\033[38;2;182;119;95m+\033[38;2;175;110;78m=\033[38;2;199;126;109m+\033[38;2;234;178;158m#\033[38;2;190;129;109m+\033[38;2;85;2;0m.\033[38;2;142;90;67m-\033[38;2;102;17;23m.\033[38;2;95;7;3m.\033[38;2;119;27;19m:\033[38;2;183;123;94m+\033[38;2;255;241;232m@\033[0m");
        $display("\033[38;2;0;0;0m          \033[38;2;21;9;5m \033[38;2;33;16;4m \033[38;2;154;136;122m+\033[38;2;198;165;144m*\033[38;2;100;60;18m:\033[38;2;255;245;219m@\033[38;2;215;186;154m#\033[38;2;203;177;138m*\033[38;2;215;188;157m#\033[38;2;138;89;51m-\033[38;2;189;150;111m*+\033[38;2;128;84;25m-\033[38;2;245;226;196m&\033[38;2;121;70;46m-\033[38;2;191;147;102m+\033[38;2;162;105;41m=\033[38;2;222;193;157m#\033[38;2;249;216;183m&\033[38;2;205;151;124m*\033[38;2;179;111;71m=\033[38;2;84;6;8m.\033[38;2;158;107;67m=\033[38;2;240;214;185m&\033[38;2;157;75;16m-\033[38;2;247;204;179m&\033[38;2;209;152;123m*\033[38;2;115;1;2m.\033[38;2;224;164;129m*\033[38;2;249;189;168m#\033[38;2;226;167;141m##\033[38;2;239;184;153m#\033[38;2;232;176;149m#\033[38;2;244;196;166m#\033[38;2;249;198;184m&\033[38;2;214;159;140m*\033[38;2;162;86;64m=\033[38;2;146;67;43m-\033[38;2;93;2;0m..\033[38;2;99;1;1m.\033[38;2;100;2;5m.\033[38;2;235;152;141m*\033[38;2;229;182;155m#\033[38;2;231;179;161m#\033[38;2;221;155;138m*\033[38;2;218;153;136m*\033[38;2;235;169;156m#\033[38;2;229;161;145m*\033[38;2;201;132;113m+\033[38;2;197;134;117m+\033[38;2;217;167;152m*\033[38;2;111;17;13m.\033[38;2;78;0;1m \033[38;2;98;25;17m.\033[38;2;119;55;40m:\033[38;2;167;118;104m+\033[38;2;153;105;91m=\033[38;2;115;51;24m:\033[38;2;112;54;30m:\033[38;2;161;119;100m=\033[38;2;105;53;34m:\033[38;2;161;124;115m+\033[38;2;62;18;10m.\033[38;2;57;2;1m \033[38;2;78;10;0m.\033[38;2;161;115;94m=\033[38;2;91;51;15m:\033[38;2;126;98;76m=\033[38;2;26;6;1m \033[38;2;28;9;8m \033[38;2;35;10;7m \033[38;2;1;2;1m    \033[38;2;3;1;2m \033[38;2;0;0;0m     \033[38;2;1;1;1m  \033[38;2;28;2;3m \033[38;2;41;1;0m \033[38;2;62;6;3m \033[38;2;79;4;1m.\033[38;2;104;21;14m.\033[38;2;99;5;5m.\033[38;2;92;4;2m.\033[38;2;96;3;0m.\033[38;2;113;11;10m.\033[38;2;160;83;63m=\033[38;2;154;86;37m-\033[38;2;138;49;0m:\033[38;2;180;106;75m=\033[38;2;181;122;89m+\033[38;2;200;136;120m+\033[38;2;221;164;142m*\033[38;2;115;27;6m.\033[38;2;80;2;1m \033[38;2;121;63;58m-\033[38;2;79;45;29m:\033[38;2;80;33;28m.\033[38;2;102;11;5m.\033[38;2;163;102;79m=\033[38;2;155;96;81m=\033[0m");
        $display("\033[38;2;0;0;0m        \033[38;2;1;1;1m  \033[38;2;22;10;2m \033[38;2;102;85;55m-\033[38;2;173;155;131m*\033[38;2;136;100;59m=\033[38;2;183;150;116m*\033[38;2;239;220;204m&\033[38;2;200;169;138m*\033[38;2;253;236;208m@\033[38;2;117;60;46m:\033[38;2;184;123;108m+\033[38;2;101;51;9m:\033[38;2;125;61;34m:\033[38;2;198;159;138m*\033[38;2;195;156;123m*\033[38;2;204;155;122m*\033[38;2;121;67;3m:\033[38;2;212;179;131m#\033[38;2;255;235;208m@\033[38;2;190;144;100m+\033[38;2;172;125;89m+\033[38;2;97;29;9m.\033[38;2;80;6;0m.\033[38;2;234;197;181m#\033[38;2;166;94;66m=\033[38;2;162;86;36m-\033[38;2;244;203;175m&\033[38;2;118;20;9m.\033[38;2;129;31;1m:\033[38;2;167;108;70m=\033[38;2;182;119;92m+\033[38;2;130;36;20m:\033[38;2;101;2;1m.\033[38;2;97;1;0m.\033[38;2;102;7;3m.\033[38;2;84;8;0m. \033[38;2;90;3;1m.\033[38;2;88;13;8m.\033[38;2;63;2;0m \033[38;2;75;4;7m. \033[38;2;55;1;1m   \033[38;2;138;49;35m:\033[38;2;217;166;144m*\033[38;2;200;128;104m+\033[38;2;220;155;136m*\033[38;2;235;174;156m#\033[38;2;228;167;146m#\033[38;2;193;131;103m+\033[38;2;180;112;92m+\033[38;2;154;88;59m=\033[38;2;134;58;14m:\033[38;2;166;108;80m=\033[38;2;174;126;109m+\033[38;2;152;102;79m=\033[38;2;85;30;22m.\033[38;2;46;2;2m \033[38;2;43;10;5m \033[38;2;37;3;2m \033[38;2;34;2;0m  \033[38;2;37;6;1m \033[38;2;41;12;7m \033[38;2;53;13;0m \033[38;2;67;3;3m \033[38;2;95;49;15m:\033[38;2;115;73;41m-\033[38;2;102;67;27m:\033[38;2;89;53;29m:\033[38;2;54;20;13m.\033[38;2;33;6;9m \033[38;2;3;0;0m   \033[38;2;1;1;1m  \033[38;2;0;0;0m    \033[38;2;1;1;1m   \033[38;2;23;3;2m \033[38;2;48;8;1m \033[38;2;73;3;3m \033[38;2;106;34;18m:\033[38;2;100;15;0m.\033[38;2;106;14;5m.\033[38;2;101;3;4m.\033[38;2;100;6;5m.\033[38;2;137;60;48m-\033[38;2;116;24;0m.\033[38;2;145;60;17m-\033[38;2;147;73;24m-\033[38;2;168;101;75m=\033[38;2;185;121;95m++\033[38;2;154;87;41m-\033[38;2;180;116;91m+\033[38;2;107;11;4m.\033[38;2;93;3;2m.\033[38;2;107;20;9m.\033[38;2;101;19;7m.\033[38;2;88;5;3m.\033[38;2;83;0;0m \033[38;2;145;65;42m-\033[0m");
        $display("\033[38;2;1;1;1m  \033[38;2;12;12;12m \033[38;2;0;0;0m      \033[38;2;6;11;2m \033[38;2;73;67;47m:\033[38;2;190;173;152m*\033[38;2;138;112;68m=\033[38;2;97;59;9m:\033[38;2;245;225;204m&\033[38;2;206;181;149m#\033[38;2;193;162;134m*\033[38;2;192;154;140m*\033[38;2;94;43;16m:\033[38;2;137;86;55m-\033[38;2;112;58;11m:\033[38;2;120;81;35m-\033[38;2;204;169;142m*\033[38;2;141;100;49m=\033[38;2;131;83;10m-\033[38;2;201;167;123m*\033[38;2;255;237;215m@\033[38;2;216;186;149m#\033[38;2;172;130;91m+\033[38;2;96;29;0m.\033[38;2;65;0;4m .\033[38;2;207;163;147m*\033[38;2;116;33;5m:\033[38;2;219;173;148m#\033[38;2;189;126;90m+\033[38;2;105;7;3m.\033[38;2;115;8;0m..\033[38;2;140;61;38m-\033[38;2;198;142;111m+\033[38;2;226;174;152m#\033[38;2;235;186;171m#\033[38;2;241;194;176m#\033[38;2;235;193;177m#\033[38;2;217;175;154m#\033[38;2;214;173;146m#\033[38;2;206;153;141m*\033[38;2;191;143;130m*\033[38;2;180;133;110m+\033[38;2;173;116;104m+=\033[38;2;134;69;40m-\033[38;2;99;9;1m.\033[38;2;127;29;10m:\033[38;2;195;129;110m+\033[38;2;177;104;72m=\033[38;2;218;147;123m*\033[38;2;233;172;151m#\033[38;2;253;205;187m&\033[38;2;221;161;147m*\033[38;2;157;81;49m-\033[38;2;126;27;3m:\033[38;2;202;140;121m*\033[38;2;168;110;97m=\033[38;2;69;1;0m  \033[38;2;58;23;19m.\033[38;2;222;215;209m&\033[38;2;85;72;68m:\033[38;2;29;0;0m \033[38;2;18;12;6m \033[38;2;28;2;2m \033[38;2;32;3;0m \033[38;2;39;11;4m \033[38;2;45;19;8m.\033[38;2;53;5;0m \033[38;2;87;20;11m.\033[38;2;117;71;38m-\033[38;2;133;92;68m-\033[38;2;87;46;6m:\033[38;2;139;110;90m=\033[38;2;51;18;5m.\033[38;2;5;0;0m   \033[38;2;1;1;1m  \033[38;2;0;0;0m     \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;22;3;2m \033[38;2;49;8;4m \033[38;2;76;2;2m \033[38;2;95;14;7m.\033[38;2;134;56;44m-\033[38;2;103;11;2m.\033[38;2;102;3;0m.\033[38;2;107;0;1m.\033[38;2;123;46;13m:\033[38;2;125;51;6m:\033[38;2;147;67;7m-\033[38;2;168;95;62m==\033[38;2;167;99;75m=\033[38;2;152;81;41m-\033[38;2;134;70;27m-\033[38;2;136;62;23m-\033[38;2;149;83;49m-\033[38;2;150;71;34m-\033[38;2;189;128;100m+\033[38;2;174;110;93m=\033[38;2;190;130;102m+\033[38;2;220;163;148m*\033[38;2;188;132;112m+\033[0m");
        $display("\033[38;2;2;2;2m \033[38;2;30;30;30m.\033[38;2;4;4;4m \033[38;2;1;1;1m \033[38;2;0;0;0m   \033[38;2;2;1;6m \033[38;2;9;6;1m \033[38;2;33;31;10m.\033[38;2;120;104;82m=\033[38;2;132;120;89m=\033[38;2;97;53;37m:\033[38;2;142;97;80m=\033[38;2;240;223;193m&\033[38;2;192;157;125m*\033[38;2;233;213;191m&\033[38;2;65;4;0m \033[38;2;148;116;93m=\033[38;2;69;8;8m.\033[38;2;104;50;9m:\033[38;2;165;128;84m+\033[38;2;130;89;42m-\033[38;2;152;111;59m=\033[38;2;196;158;112m*\033[38;2;232;212;175m&\033[38;2;219;194;162m#\033[38;2;167;108;65m=\033[38;2;97;24;17m.\033[38;2;62;2;6m \033[38;2;56;1;0m \033[38;2;210;169;155m*\033[38;2;160;113;66m=\033[38;2;106;23;12m.\033[38;2;247;203;180m&\033[38;2;128;42;1m:\033[38;2;92;1;0m.\033[38;2;104;7;2m.\033[38;2;178;117;97m+\033[38;2;201;152;130m**\033[38;2;196;130;111m+\033[38;2;224;158;134m*\033[38;2;176;106;76m=\033[38;2;164;98;65m=\033[38;2;189;130;102m+\033[38;2;141;79;55m-\033[38;2;125;46;27m:\033[38;2;88;13;13m..\033[38;2;69;1;2m \033[38;2;142;71;58m-\033[38;2;191;151;135m*\033[38;2;190;138;121m+\033[38;2;103;8;0m.\033[38;2;136;44;19m:\033[38;2;169;87;62m=\033[38;2;221;165;142m*\033[38;2;237;178;159m#\033[38;2;246;183;162m#\033[38;2;244;186;170m#\033[38;2;150;66;18m-\033[38;2;121;15;2m.\033[38;2;122;30;17m:\033[38;2;74;8;5m.\033[38;2;69;0;0m \033[38;2;122;62;36m:\033[38;2;89;27;10m.\033[38;2;46;4;1m \033[38;2;50;9;9m \033[38;2;43;7;0m  \033[38;2;68;8;1m \033[38;2;136;96;74m=\033[38;2;193;159;135m*\033[38;2;50;3;1m \033[38;2;48;2;5m \033[38;2;54;0;0m \033[38;2;70;9;1m.\033[38;2;133;88;40m-\033[38;2;147;106;82m=\033[38;2;64;5;1m \033[38;2;70;36;31m.\033[38;2;21;4;3m \033[38;2;4;0;1m           \033[38;2;34;1;2m \033[38;2;58;8;5m \033[38;2;78;6;0m.\033[38;2;103;29;18m.\033[38;2;124;52;24m:\033[38;2;114;39;8m:.\033[38;2;121;34;5m::\033[38;2;107;4;0m.\033[38;2;147;66;24m-\033[38;2;179;114;78m=\033[38;2;147;73;36m-\033[38;2;137;54;9m:\033[38;2;118;34;8m:\033[38;2;123;50;6m:\033[38;2;146;63;31m-\033[38;2;126;49;9m:\033[38;2;142;54;32m-\033[38;2;174;87;72m=\033[38;2;184;108;92m=\033[38;2;123;36;26m:\033[38;2;106;5;0m.\033[38;2;143;68;47m-\033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m   \033[38;2;2;6;1m \033[38;2;5;18;3m \033[38;2;29;32;14m.\033[38;2;55;43;20m.\033[38;2;195;176;161m*\033[38;2;171;151;124m+\033[38;2;60;2;0m \033[38;2;187;162;131m*\033[38;2;197;167;134m*\033[38;2;183;156;130m*\033[38;2;67;16;5m.\033[38;2;114;71;52m-\033[38;2;59;10;2m .\033[38;2;87;30;4m.\033[38;2;127;90;39m-\033[38;2;139;96;46m-\033[38;2;160;117;76m=\033[38;2;214;182;153m#\033[38;2;255;241;208m@\033[38;2;151;109;53m=\033[38;2;77;7;3m.\033[38;2;105;51;36m:\033[38;2;54;3;2m \033[38;2;83;11;3m.\033[38;2;198;158;131m*\033[38;2;96;8;1m.\033[38;2;147;93;56m=\033[38;2;181;124;88m+\033[38;2;101;8;1m.\033[38;2;132;50;20m:\033[38;2;111;20;0m.\033[38;2;185;116;94m+\033[38;2;182;118;95m+\033[38;2;178;103;76m=\033[38;2;140;68;50m-\033[38;2;148;82;65m-\033[38;2;93;8;5m.\033[38;2;57;3;1m \033[38;2;51;20;13m.\033[38;2;32;5;0m \033[38;2;22;10;4m \033[38;2;72;55;50m:\033[38;2;52;17;10m.\033[38;2;51;3;4m \033[38;2;49;20;5m.\033[38;2;58;8;4m \033[38;2;102;11;6m.\033[38;2;115;13;10m.\033[38;2;124;17;9m.\033[38;2;165;89;53m=\033[38;2;202;119;98m+\033[38;2;190;112;73m+\033[38;2;233;159;135m*\033[38;2;203;134;113m+\033[38;2;223;159;144m*\033[38;2;154;61;40m-\033[38;2;122;25;3m.\033[38;2;145;56;37m-\033[38;2;182;120;105m+\033[38;2;151;84;43m-\033[38;2;162;98;71m=\033[38;2;142;79;57m-\033[38;2;149;90;68m=\033[38;2;155;99;83m==\033[38;2;149;89;62m=\033[38;2;175;110;83m=\033[38;2;172;126;98m+\033[38;2;153;105;77m=\033[38;2;63;2;1m \033[38;2;54;0;0m \033[38;2;65;8;4m \033[38;2;105;55;26m:\033[38;2;135;97;72m=\033[38;2;62;14;5m.\033[38;2;42;15;3m \033[38;2;23;2;0m \033[38;2;10;0;3m \033[38;2;0;2;1m            \033[38;2;88;19;10m.\033[38;2;113;47;26m:\033[38;2;133;61;32m-\033[38;2;119;41;9m:\033[38;2;139;61;37m-\033[38;2;144;67;35m-\033[38;2;145;61;33m-\033[38;2;129;54;1m:\033[38;2;154;80;40m-\033[38;2;143;67;38m-\033[38;2;139;70;46m-\033[38;2;92;2;0m..\033[38;2;89;9;3m.\033[38;2;86;5;2m.\033[38;2;113;45;37m:\033[38;2;103;29;31m.\033[38;2;97;25;33m.\033[38;2;109;40;48m:\033[38;2;70;9;8m.\033[38;2;69;2;1m \033[38;2;126;55;55m:\033[0m");
        $display("\033[38;2;0;0;0m       \033[38;2;13;25;8m \033[38;2;25;10;1m \033[38;2;168;149;121m+\033[38;2;86;59;19m:\033[38;2;88;50;10m:\033[38;2;74;13;14m.\033[38;2;215;190;174m#\033[38;2;160;131;90m+\033[38;2;141;107;81m=\033[38;2;51;2;0m \033[38;2;88;45;34m:\033[38;2;44;2;1m \033[38;2;88;34;17m.\033[38;2;84;27;3m.\033[38;2;106;52;12m:\033[38;2;116;73;18m-\033[38;2;184;145;116m+\033[38;2;254;233;210m@\033[38;2;170;132;97m+\033[38;2;63;1;5m \033[38;2;116;58;51m:\033[38;2;73;18;9m.\033[38;2;68;2;2m \033[38;2;85;30;17m.\033[38;2;155;95;77m=\033[38;2;108;24;11m.\033[38;2;158;90;70m=\033[38;2;137;70;15m-\033[38;2;142;75;17m-\033[38;2;129;41;8m:\033[38;2;136;55;32m:\033[38;2;161;98;71m=\033[38;2;155;97;73m=\033[38;2;140;77;63m-\033[38;2;63;6;5m \033[38;2;60;21;12m.\033[38;2;35;2;2m  \033[38;2;40;10;9m \033[38;2;49;34;27m.\033[38;2;43;6;6m \033[38;2;203;174;166m#\033[38;2;58;25;16m.\033[38;2;46;5;1m \033[38;2;92;31;25m.\033[38;2;179;140;112m+\033[38;2;125;60;27m:\033[38;2;153;85;49m-\033[38;2;161;94;69m=\033[38;2;193;114;81m+\033[38;2;186;99;68m=\033[38;2;191;119;92m+\033[38;2;203;130;108m++\033[38;2;202;128;114m+\033[38;2;231;157;150m*\033[38;2;165;67;55m-\033[38;2;127;6;0m.\033[38;2;160;80;59m-\033[38;2;195;124;110m+\033[38;2;200;132;109m+\033[38;2;207;138;123m*\033[38;2;181;109;95m=\033[38;2;180;110;99m+\033[38;2;185;117;104m+\033[38;2;195;128;112m+\033[38;2;177;110;91m=\033[38;2;169;105;76m=\033[38;2;174;118;96m+\033[38;2;153;97;81m=\033[38;2;68;3;0m \033[38;2;65;0;1m \033[38;2;72;8;3m.\033[38;2;127;85;60m-\033[38;2;99;47;34m:\033[38;2;47;12;5m \033[38;2;32;1;0m \033[38;2;24;6;4m \033[38;2;1;1;1m \033[38;2;0;0;0m          \033[38;2;46;1;1m \033[38;2;92;35;28m.\033[38;2;99;28;4m.\033[38;2;115;42;9m:\033[38;2;137;68;38m-\033[38;2;136;66;18m-\033[38;2;152;81;52m-\033[38;2;166;94;64m=\033[38;2;160;101;62m==\033[38;2;149;81;48m-\033[38;2;124;43;31m:\033[38;2;62;14;9m.\033[38;2;63;25;19m.\033[38;2;50;10;3m \033[38;2;59;9;11m \033[38;2;50;6;2m  \033[38;2;49;4;6m \033[38;2;43;2;1m \033[38;2;46;1;0m \033[38;2;48;2;2m \033[38;2;49;5;4m \033[0m");
        $display("\033[38;2;0;0;0m    \033[38;2;1;1;1m \033[38;2;6;6;4m \033[38;2;0;0;2m \033[38;2;36;37;17m.\033[38;2;118;98;81m-\033[38;2;146;130;104m+\033[38;2;87;47;19m:\033[38;2;60;4;1m \033[38;2;171;139;114m+\033[38;2;214;182;158m#\033[38;2;175;143;103m+\033[38;2;62;4;1m \033[38;2;57;5;3m \033[38;2;55;0;1m  \033[38;2;86;33;14m.\033[38;2;89;31;4m.\033[38;2;100;43;0m:\033[38;2;134;99;35m-\033[38;2;227;192;170m#\033[38;2;238;202;178m&\033[38;2;61;3;1m \033[38;2;109;64;54m:\033[38;2;56;3;1m \033[38;2;71;2;2m \033[38;2;91;19;11m.\033[38;2;170;126;91m+\033[38;2;102;17;3m.\033[38;2;97;9;0m.\033[38;2;180;123;91m+\033[38;2;167;102;69m=\033[38;2;150;77;42m-\033[38;2;145;69;34m-\033[38;2;109;15;5m.\033[38;2;155;71;47m-\033[38;2;189;124;101m+\033[38;2;139;66;48m-\033[38;2;124;56;45m:\033[38;2;128;62;57m-\033[38;2;74;7;1m.\033[38;2;81;19;8m.\033[38;2;73;2;0m \033[38;2;117;35;15m:\033[38;2;159;97;76m=\033[38;2;172;116;102m+\033[38;2;178;118;114m+\033[38;2;195;136;123m+\033[38;2;176;102;82m=\033[38;2;186;109;87m+\033[38;2;175;93;73m=\033[38;2;194;122;105m+\033[38;2;188;111;94m+\033[38;2;165;81;35m-\033[38;2;192;114;84m+\033[38;2;210;136;112m+\033[38;2;213;142;123m*\033[38;2;208;137;113m+\033[38;2;211;136;116m*\033[38;2;229;162;145m*\033[38;2;200;134;118m+\033[38;2;180;90;63m=\033[38;2;123;5;0m.\033[38;2;169;96;70m=\033[38;2;198;118;98m+\033[38;2;205;135;116m+\033[38;2;225;153;138m*\033[38;2;214;147;131m*\033[38;2;213;141;127m*\033[38;2;209;140;124m*\033[38;2;185;119;97m+\033[38;2;180;108;93m=\033[38;2;166;99;73m=\033[38;2;140;79;53m-\033[38;2;88;14;3m.\033[38;2;59;0;1m \033[38;2;65;1;0m \033[38;2;112;65;42m:\033[38;2;151;120;94m=\033[38;2;48;0;1m \033[38;2;31;10;3m \033[38;2;29;3;4m \033[38;2;8;0;1m  \033[38;2;3;1;2m \033[38;2;1;0;0m       \033[38;2;26;1;2m \033[38;2;43;8;6m .\033[38;2;106;41;24m:\033[38;2;112;44;8m:\033[38;2;133;67;32m-\033[38;2;124;50;2m:\033[38;2;137;58;4m:\033[38;2;142;66;10m-\033[38;2;135;62;8m-\033[38;2;141;61;25m-\033[38;2;119;47;3m:\033[38;2;108;31;6m.\033[38;2;94;8;0m.\033[38;2;89;13;13m.\033[38;2;139;83;74m-\033[38;2;250;234;224m@\033[38;2;254;248;245m@\033[38;2;247;251;249m@\033[38;2;215;172;172m#\033[38;2;196;145;146m*\033[38;2;177;127;128m+\033[38;2;80;34;34m.\033[38;2;114;78;83m-\033[0m");
        $display("\033[38;2;0;0;0m      \033[38;2;14;16;8m \033[38;2;24;25;13m \033[38;2;126;117;82m=\033[38;2;106;76;41m-\033[38;2;70;22;10m.\033[38;2;129;97;50m-\033[38;2;162;138;110m+\033[38;2;170;140;105m+\033[38;2;66;8;2m  \033[38;2;76;9;1m.\033[38;2;53;2;0m \033[38;2;51;0;1m \033[38;2;74;19;11m.\033[38;2;64;1;1m \033[38;2;99;42;13m:\033[38;2;180;152;123m*\033[38;2;203;174;143m*\033[38;2;62;5;2m \033[38;2;51;2;0m \033[38;2;92;42;25m:\033[38;2;47;4;2m  \033[38;2;113;52;47m:\033[38;2;95;26;13m.\033[38;2;103;18;3m.\033[38;2;153;93;42m=\033[38;2;143;61;8m-\033[38;2;131;48;17m:\033[38;2;154;80;53m-\033[38;2;152;76;41m-\033[38;2;123;38;12m:\033[38;2;165;102;73m=\033[38;2;180;114;80m+\033[38;2;217;155;137m*\033[38;2;210;143;127m*\033[38;2;209;140;121m*\033[38;2;181;116;90m+\033[38;2;192;134;109m+\033[38;2;178;115;98m+\033[38;2;216;155;146m*\033[38;2;207;134;109m+\033[38;2;210;138;113m*\033[38;2;197;125;100m+\033[38;2;201;121;104m++\033[38;2;195;112;96m+\033[38;2;180;101;86m=\033[38;2;220;143;133m*\033[38;2;221;139;131m*\033[38;2;211;138;117m*\033[38;2;226;159;140m**\033[38;2;206;131;108m+\033[38;2;207;130;110m+\033[38;2;220;146;134m*\033[38;2;229;156;147m*\033[38;2;224;155;132m*\033[38;2;194;122;107m+\033[38;2;163;74;40m--\033[38;2;210;141;120m*\033[38;2;206;139;123m*\033[38;2;214;145;130m*\033[38;2;227;154;143m*\033[38;2;199;128;111m+\033[38;2;210;136;125m*\033[38;2;194;121;106m++\033[38;2;198;131;115m+\033[38;2;151;81;63m-\033[38;2;117;53;18m:\033[38;2;67;0;0m  \033[38;2;81;23;4m.\033[38;2;117;84;53m-\033[38;2;88;50;43m:\033[38;2;36;4;5m \033[38;2;28;0;0m  \033[38;2;26;2;8m \033[38;2;13;1;6m \033[38;2;2;0;1m        \033[38;2;40;2;0m \033[38;2;50;4;3m \033[38;2;115;54;42m:\033[38;2;103;32;6m.\033[38;2;125;61;26m:\033[38;2;139;71;32m-\033[38;2;140;69;40m-\033[38;2;147;75;39m--\033[38;2;121;50;6m:\033[38;2;134;70;21m-\033[38;2;96;11;14m.\033[38;2;121;46;23m:\033[38;2;228;178;160m#\033[38;2;254;219;204m&\033[38;2;243;205;188m&\033[38;2;197;124;96m+\033[38;2;169;64;46m-\033[38;2;113;8;6m.\033[38;2;98;3;2m.\033[38;2;141;67;56m-\033[38;2;205;151;139m*\033[38;2;224;199;190m#\033[0m");
        $display("\033[38;2;0;0;0m    \033[38;2;2;2;1m \033[38;2;21;21;13m \033[38;2;44;42;23m.\033[38;2;79;73;40m:\033[38;2;116;94;63m-\033[38;2;84;49;4m::\033[38;2;128;98;59m-\033[38;2;137;110;80m=\033[38;2;125;86;59m-\033[38;2;67;2;4m \033[38;2;97;52;34m:\033[38;2;45;1;0m  \033[38;2;49;3;1m   \033[38;2;155;117;80m=\033[38;2;187;152;122m*\033[38;2;85;36;22m.\033[38;2;71;29;26m.\033[38;2;96;58;42m:\033[38;2;52;14;5m \033[38;2;53;21;4m.\033[38;2;109;51;37m:\033[38;2;97;39;19m:\033[38;2;83;7;4m.\033[38;2;113;36;19m:\033[38;2;136;61;21m-\033[38;2;134;54;6m:\033[38;2;138;55;12m:\033[38;2;142;66;15m-\033[38;2;153;76;34m-\033[38;2;173;104;64m=\033[38;2;215;153;132m*\033[38;2;180;112;81m=\033[38;2;207;142;111m*\033[38;2;204;138;115m+\033[38;2;197;132;111m+\033[38;2;238;174;159m#\033[38;2;233;169;151m#\033[38;2;218;150;131m*\033[38;2;229;151;138m*\033[38;2;216;144;132m*\033[38;2;220;143;131m*\033[38;2;214;133;121m*\033[38;2;209;129;118m+\033[38;2;214;137;122m*\033[38;2;240;165;152m#\033[38;2;239;169;161m#\033[38;2;242;170;160m#\033[38;2;202;109;96m+\033[38;2;215;143;121m**\033[38;2;209;131;106m+\033[38;2;174;94;61m=\033[38;2;192;114;92m+\033[38;2;211;136;118m*\033[38;2;227;155;145m*\033[38;2;230;168;161m#\033[38;2;218;151;132m*\033[38;2;171;92;70m=\033[38;2;168;70;54m-\033[38;2;164;61;40m-\033[38;2;189;112;89m+\033[38;2;212;139;122m*\033[38;2;222;160;145m*\033[38;2;218;148;135m*\033[38;2;220;149;137m*\033[38;2;207;135;123m+\033[38;2;193;124;107m+\033[38;2;192;123;108m+\033[38;2;154;81;48m-\033[38;2;130;75;45m-\033[38;2;95;24;13m.\033[38;2;64;0;1m \033[38;2;71;13;2m.\033[38;2;84;38;12m.\033[38;2;103;58;51m:\033[38;2;31;13;3m   \033[38;2;2;2;2m  \033[38;2;0;1;0m     \033[38;2;2;2;2m \033[38;2;10;0;1m  \033[38;2;30;2;0m \033[38;2;36;0;2m \033[38;2;69;15;4m.\033[38;2;81;8;5m.\033[38;2;112;43;14m:\033[38;2;115;44;6m:\033[38;2;134;57;16m:\033[38;2;141;69;29m-\033[38;2;127;51;7m:\033[38;2;112;21;6m.\033[38;2;199;141;123m*\033[38;2;218;189;171m#\033[38;2;255;252;241m@\033[38;2;254;227;203m&\033[38;2;250;214;188m&\033[38;2;253;217;197m&\033[38;2;255;208;190m&&\033[38;2;248;190;173m#\033[38;2;243;192;175m#\033[38;2;238;213;189m&\033[38;2;240;192;175m#\033[38;2;233;184;173m#\033[0m");
        $display("\033[38;2;5;3;4m \033[38;2;85;81;82m-\033[38;2;137;131;133m+\033[38;2;248;247;242m@\033[38;2;238;234;223m@\033[38;2;227;215;201m&\033[38;2;196;178;164m#\033[38;2;113;88;50m-\033[38;2;101;71;17m:\033[38;2;98;60;1m:\033[38;2;104;63;15m:\033[38;2;120;86;26m-\033[38;2;142;106;70m=\033[38;2;81;20;0m. \033[38;2;109;70;52m-\033[38;2;56;5;3m \033[38;2;53;3;2m \033[38;2;42;0;3m  \033[38;2;85;32;11m.\033[38;2;169;134;109m+\033[38;2;141;98;71m=\033[38;2;53;0;1m \033[38;2;52;1;0m \033[38;2;118;76;57m-\033[38;2;50;8;2m \033[38;2;46;11;0m \033[38;2;127;75;62m-\033[38;2;113;52;29m:\033[38;2;82;0;0m \033[38;2;125;56;21m:\033[38;2;119;47;4m:\033[38;2;130;50;0m:\033[38;2;138;40;5m:\033[38;2;172;107;78m=\033[38;2;189;117;93m++\033[38;2;187;114;91m+\033[38;2;197;125;104m+\033[38;2;192;114;94m+\033[38;2;212;136;111m*\033[38;2;219;148;124m*\033[38;2;222;151;130m*\033[38;2;226;154;138m*\033[38;2;235;162;146m#\033[38;2;228;159;144m*\033[38;2;224;156;145m*\033[38;2;237;162;151m#\033[38;2;239;169;157m#\033[38;2;248;171;161m#\033[38;2;238;162;150m#\033[38;2;241;173;158m#\033[38;2;250;177;166m#\033[38;2;242;169;162m#\033[38;2;208;133;120m+\033[38;2;187;106;77m=\033[38;2;158;67;25m-\033[38;2;172;80;46m=\033[38;2;159;58;28m-\033[38;2;178;75;39m-\033[38;2;209;123;109m+\033[38;2;215;146;131m*\033[38;2;237;166;157m#\033[38;2;250;221;217m&&\033[38;2;217;156;140m*\033[38;2;174;106;74m=\033[38;2;136;43;7m:\033[38;2;171;88;64m=\033[38;2;193;116;106m+\033[38;2;197;129;110m+\033[38;2;198;121;103m+\033[38;2;193;115;97m+\033[38;2;177;105;85m=\033[38;2;167;96;76m=\033[38;2;164;91;73m=\033[38;2;119;71;35m-\033[38;2;92;33;13m.\033[38;2;58;0;3m \033[38;2;68;15;7m.\033[38;2;63;7;1m \033[38;2;128;99;87m=\033[38;2;44;23;8m.\033[38;2;29;2;3m  \033[38;2;7;1;1m   \033[38;2;0;0;0m    \033[38;2;2;2;2m  \033[38;2;8;0;0m  \033[38;2;34;1;2m \033[38;2;41;5;0m   \033[38;2;78;2;1m \033[38;2;147;71;45m-\033[38;2;191;143;108m+\033[38;2;234;198;169m#\033[38;2;255;246;237m@\033[38;2;253;250;240m@\033[38;2;251;228;216m@&\033[38;2;254;194;173m&&&&\033[38;2;255;202;188m&\033[38;2;254;198;178m&\033[38;2;240;168;148m#\033[38;2;199;132;105m+\033[38;2;211;145;119m*\033[38;2;233;182;160m#\033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;236;234;235m@\033[38;2;240;218;224m&\033[38;2;210;176;176m#\033[38;2;198;164;156m**\033[38;2;188;148;126m*\033[38;2;140;91;61m-\033[38;2;95;42;0m:.\033[38;2;96;47;5m:\033[38;2;149;109;80m=\033[38;2;142;100;59m=\033[38;2;75;6;2m.\033[38;2;61;2;3m \033[38;2;135;91;71m-\033[38;2;53;2;3m \033[38;2;55;3;0m \033[38;2;53;1;1m  \033[38;2;116;67;32m-\033[38;2;131;95;70m-\033[38;2;75;23;4m.\033[38;2;51;1;2m \033[38;2;68;14;14m.\033[38;2;94;55;37m:\033[38;2;40;13;1m \033[38;2;58;25;6m.\033[38;2;139;96;88m=\033[38;2;96;38;7m:\033[38;2;99;16;5m.\033[38;2;125;48;18m:\033[38;2;100;7;0m.:\033[38;2;136;55;9m:\033[38;2;172;92;67m===\033[38;2;171;95;64m=\033[38;2;165;90;59m=\033[38;2;176;99;71m=\033[38;2;201;124;101m+\033[38;2;191;120;94m+\033[38;2;199;128;102m+\033[38;2;200;124;100m+\033[38;2;208;131;111m+\033[38;2;223;150;143m*\033[38;2;245;180;168m#\033[38;2;241;165;156m#\033[38;2;250;181;170m#\033[38;2;249;186;171m#\033[38;2;244;173;160m##\033[38;2;249;181;172m#\033[38;2;210;129;112m+\033[38;2;190;97;83m=\033[38;2;163;68;42m-\033[38;2;164;69;52m-\033[38;2;195;131;112m+\033[38;2;219;161;153m*\033[38;2;193;125;111m+\033[38;2;126;35;26m:\033[38;2;129;24;15m:\033[38;2;178;106;87m=\033[38;2;192;104;84m=\033[38;2;178;88;65m=\033[38;2;186;102;82m=\033[38;2;164;77;51m-\033[38;2;116;0;0m.\033[38;2;178;101;85m=\033[38;2;203;128;114m+\033[38;2;177;97;81m=\033[38;2;179;90;77m=\033[38;2;185;106;89m=\033[38;2;187;115;95m+\033[38;2;167;96;75m=\033[38;2;136;66;39m-\033[38;2;100;30;6m.\033[38;2;97;41;21m:\033[38;2;70;1;3m \033[38;2;62;2;2m \033[38;2;68;9;3m.\033[38;2;108;72;62m-\033[38;2;40;14;3m \033[38;2;23;1;2m \033[38;2;30;4;3m  \033[38;2;9;2;2m \033[38;2;5;0;4m    \033[38;2;1;1;1m \033[38;2;2;2;2m   \033[38;2;44;21;17m.\033[38;2;48;29;15m.\033[38;2;90;52;44m:\033[38;2;149;105;91m=\033[38;2;211;181;158m#\033[38;2;230;205;190m&\033[38;2;251;238;226m@\033[38;2;254;246;239m@\033[38;2;255;242;223m@\033[38;2;249;218;207m&\033[38;2;230;178;157m#\033[38;2;236;175;150m#\033[38;2;243;176;155m##\033[38;2;251;182;159m#\033[38;2;252;188;165m#\033[38;2;250;192;170m##\033[38;2;249;188;163m#\033[38;2;242;175;150m#\033[38;2;233;162;138m*\033[38;2;231;165;139m#\033[38;2;247;197;171m&\033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;198;187;187m#\033[38;2;216;178;169m#\033[38;2;195;157;137m*\033[38;2;174;122;108m+\033[38;2;193;152;131m*\033[38;2;159;119;97m==\033[38;2;94;44;4m:\033[38;2;85;32;1m.\033[38;2;125;77;28m-\033[38;2;131;91;50m-\033[38;2;128;92;49m-\033[38;2;81;23;1m. \033[38;2;125;81;48m-\033[38;2;69;8;3m.\033[38;2;76;5;2m.\033[38;2;64;0;1m \033[38;2;63;1;2m \033[38;2;130;85;48m-\033[38;2;146;106;77m=\033[38;2;82;17;2m.\033[38;2;61;1;1m  \033[38;2;103;54;24m:\033[38;2;61;2;0m \033[38;2;50;0;2m \033[38;2;124;77;58m-\033[38;2;98;35;12m.\033[38;2;86;0;0m.\033[38;2;96;14;3m.\033[38;2;87;2;4m.\033[38;2;104;27;6m.\033[38;2;142;73;21m-\033[38;2;145;67;23m-\033[38;2;150;62;24m-\033[38;2;155;78;56m-\033[38;2;176;109;81m=\033[38;2;174;107;76m=\033[38;2;170;90;63m=\033[38;2;179;95;66m=\033[38;2;180;102;82m=\033[38;2;183;98;76m=\033[38;2;181;96;75m=\033[38;2;190;105;76m=\033[38;2;204;126;104m+\033[38;2;218;146;128m*\033[38;2;221;152;136m***\033[38;2;231;160;144m**\033[38;2;228;156;140m*\033[38;2;178;80;47m=\033[38;2;217;138;125m*\033[38;2;123;10;2m.\033[38;2;114;4;1m.\033[38;2;125;12;13m.\033[38;2;93;0;4m.\033[38;2;95;36;35m:\033[38;2;70;14;13m.\033[38;2;102;0;0m.\033[38;2;115;3;1m.\033[38;2;130;13;10m.\033[38;2;110;3;1m..\033[38;2;152;94;68m=\033[38;2;177;113;96m+\033[38;2;163;92;73m=\033[38;2;177;111;85m=\033[38;2;192;133;117m+\033[38;2;160;76;48m-\033[38;2;185;107;95m=\033[38;2;175;109;83m=\033[38;2;163;96;70m=\033[38;2;130;56;16m:\033[38;2;107;45;9m:\033[38;2;77;13;1m.\033[38;2;70;12;8m.\033[38;2;55;6;3m .\033[38;2;66;32;17m.\033[38;2;27;12;5m \033[38;2;22;2;1m  \033[38;2;34;0;0m \033[38;2;28;2;3m  \033[38;2;2;0;1m    \033[38;2;3;4;4m \033[38;2;81;66;66m:\033[38;2;64;34;36m.\033[38;2;230;218;219m&\033[38;2;251;252;251m@\033[38;2;254;244;249m@\033[38;2;252;251;251m@\033[38;2;253;246;249m@@\033[38;2;252;251;233m@\033[38;2;255;220;205m&\033[38;2;251;198;167m&#&\033[38;2;253;193;165m&\033[38;2;249;185;157m#\033[38;2;241;177;149m#\033[38;2;238;174;146m##\033[38;2;234;173;145m#\033[38;2;240;179;151m#\033[38;2;247;189;159m#\033[38;2;242;178;151m#\033[38;2;237;172;146m#\033[38;2;251;186;166m#\033[38;2;241;194;171m#\033[0m");
        $display("\033[38;2;0;2;1m \033[38;2;178;163;160m*\033[38;2;182;142;131m+\033[38;2;158;112;92m=\033[38;2;147;96;71m=\033[38;2;167;123;89m+\033[38;2;134;88;50m-\033[38;2;153;107;82m=\033[38;2;98;37;10m:\033[38;2;92;38;4m.\033[38;2;119;73;29m-\033[38;2;115;74;17m-\033[38;2;130;89;46m-\033[38;2;94;35;12m.\033[38;2;103;49;4m:\033[38;2;153;119;75m=\033[38;2;117;62;6m:\033[38;2;119;76;21m-\033[38;2;101;41;7m:\033[38;2;92;29;9m.\033[38;2;128;76;25m-\033[38;2;141;97;61m=\033[38;2;98;40;9m:\033[38;2;84;18;5m.\033[38;2;79;3;4m.\033[38;2;126;75;45m-\033[38;2;86;16;2m. \033[38;2;72;3;1m \033[38;2;176;122;90m+\033[38;2;121;55;11m:\033[38;2;124;59;18m:\033[38;2;119;31;8m:\033[38;2;133;55;34m:\033[38;2;159;95;53m=\033[38;2;157;84;51m-\033[38;2;163;85;46m=\033[38;2;146;71;32m-\033[38;2;161;90;57m===\033[38;2;167;86;59m=\033[38;2;175;90;69m=\033[38;2;178;95;71m=\033[38;2;169;83;50m=\033[38;2;173;88;63m=\033[38;2;177;92;71m=\033[38;2;195;113;92m+\033[38;2;202;124;104m+\033[38;2;203;127;108m+\033[38;2;204;126;105m+\033[38;2;196;117;95m++\033[38;2;199;113;91m+\033[38;2;161;61;12m-\033[38;2;217;142;125m*\033[38;2;228;146;135m*\033[38;2;135;46;29m:\033[38;2;198;120;106m+\033[38;2;223;147;141m*\033[38;2;242;179;169m#\033[38;2;241;187;175m#\033[38;2;250;216;200m&\033[38;2;200;129;106m++\033[38;2;242;196;181m&\033[38;2;229;181;170m#\033[38;2;196;129;113m+\033[38;2;140;61;30m-:\033[38;2;152;75;45m-\033[38;2;147;54;29m-\033[38;2;215;152;141m*\033[38;2;183;122;101m+=\033[38;2;141;70;36m-\033[38;2;120;45;5m:\033[38;2;124;75;42m-\033[38;2;86;27;9m.\033[38;2;64;9;8m \033[38;2;45;13;5m \033[38;2;74;44;24m.\033[38;2;70;40;27m.\033[38;2;36;12;9m \033[38;2;26;5;2m \033[38;2;32;0;3m \033[38;2;31;2;4m \033[38;2;30;0;2m \033[38;2;6;2;0m \033[38;2;23;6;5m \033[38;2;24;8;7m \033[38;2;73;59;59m:\033[38;2;96;75;81m-\033[38;2;204;194;193m#\033[38;2;254;251;250m@\033[38;2;255;253;255m@@@\033[38;2;254;236;244m@\033[38;2;253;233;233m@@\033[38;2;250;200;190m&&\033[38;2;252;204;182m&\033[38;2;254;217;190m&&\033[38;2;251;220;202m&\033[38;2;254;205;183m&\033[38;2;249;183;157m#\033[38;2;238;174;146m###\033[38;2;230;165;137m*\033[38;2;239;175;147m#\033[38;2;250;189;162m#\033[38;2;252;188;166m#\033[38;2;254;196;170m&\033[38;2;247;181;157m#\033[38;2;248;196;173m&\033[0m");
        $display("\033[38;2;2;3;5m \033[38;2;97;73;67m-\033[38;2;116;53;36m:\033[38;2;91;9;0m..\033[38;2;119;53;23m:\033[38;2;121;63;41m-\033[38;2;143;92;63m=\033[38;2;113;58;12m:\033[38;2;72;0;1m \033[38;2;93;38;2m.\033[38;2;125;83;42m-\033[38;2;117;71;19m-\033[38;2;98;33;7m.\033[38;2;123;65;15m:\033[38;2;206;173;142m*\033[38;2;155;116;58m=\033[38;2;152;104;56m=\033[38;2;88;13;0m.\033[38;2;89;21;8m.\033[38;2;109;62;3m:\033[38;2;158;117;82m=\033[38;2;125;84;29m-\033[38;2;107;45;0m:\033[38;2;124;63;13m:\033[38;2;170;121;84m+\033[38;2;117;53;8m:\033[38;2;100;27;2m.\033[38;2;114;44;8m:\033[38;2;247;213;199m&\033[38;2;116;43;10m:\033[38;2;152;95;57m=\033[38;2;135;58;11m:\033[38;2;132;53;18m:\033[38;2;158;87;54m=\033[38;2;159;86;47m-\033[38;2;157;82;52m--\033[38;2;166;96;65m==\033[38;2;177;97;70m===\033[38;2;181;103;84m=\033[38;2;154;65;27m-\033[38;2;179;100;77m=\033[38;2;175;91;68m==\033[38;2;180;97;71m=\033[38;2;188;101;81m=\033[38;2;186;106;83m=\033[38;2;194;111;90m+\033[38;2;177;96;76m==\033[38;2;201;120;101m+\033[38;2;213;134;119m*\033[38;2;218;144;135m*\033[38;2;192;105;84m=\033[38;2;238;172;163m#\033[38;2;202;124;109m+\033[38;2;205;132;111m+\033[38;2;222;149;134m*\033[38;2;198;127;115m+\033[38;2;184;102;79m=\033[38;2;204;126;114m+\033[38;2;208;140;117m*\033[38;2;163;67;41m-\033[38;2;142;46;10m:\033[38;2;123;16;0m.\033[38;2;130;39;20m::\033[38;2;115;19;15m.\033[38;2;92;1;0m.\033[38;2;137;59;32m-\033[38;2;157;103;76m=\033[38;2;132;70;25m-\033[38;2;116;54;4m:\033[38;2;122;72;40m-\033[38;2;85;23;8m.\033[38;2;55;3;2m \033[38;2;43;1;0m \033[38;2;73;38;26m.\033[38;2;32;9;2m \033[38;2;36;1;1m    \033[38;2;35;0;4m \033[38;2;48;14;12m \033[38;2;78;59;48m:\033[38;2;197;178;177m#\033[38;2;254;253;250m@@@@\033[38;2;255;251;255m@\033[38;2;252;239;251m@\033[38;2;253;240;255m@@\033[38;2;234;188;181m#\033[38;2;241;176;162m#\033[38;2;238;170;153m#\033[38;2;242;182;150m#\033[38;2;230;158;129m*\033[38;2;255;202;177m&\033[38;2;248;197;171m&\033[38;2;251;202;178m&\033[38;2;244;182;157m#\033[38;2;243;176;150m#\033[38;2;253;192;164m#\033[38;2;240;175;147m#\033[38;2;230;166;138m#*\033[38;2;244;184;157m#\033[38;2;250;191;163m#\033[38;2;254;193;173m&\033[38;2;255;199;176m&\033[38;2;254;202;175m&&\033[0m");
        $display("\033[38;2;1;1;3m \033[38;2;108;83;79m-\033[38;2;107;47;31m:\033[38;2;106;35;2m:\033[38;2;110;46;5m:\033[38;2;115;51;9m:\033[38;2;99;39;4m:\033[38;2;112;56;13m:\033[38;2;105;46;1m:\033[38;2;116;65;35m:\033[38;2;94;26;8m.\033[38;2;116;64;21m:\033[38;2;123;81;20m-\033[38;2;96;20;5m.\033[38;2;137;90;45m-\033[38;2;215;184;154m#\033[38;2;183;147;105m+\033[38;2;147;96;51m=\033[38;2;98;39;6m:\033[38;2;60;2;1m \033[38;2;105;61;12m:\033[38;2;133;76;23m-\033[38;2;126;77;12m-\033[38;2;131;75;6m-\033[38;2;185;132;87m+\033[38;2;172;122;80m+\033[38;2;145;86;48m-\033[38;2;74;4;3m \033[38;2;83;1;0m \033[38;2;124;60;23m:\033[38;2;228;192;167m#\033[38;2;82;4;11m.\033[38;2;114;34;9m:\033[38;2;109;20;0m.\033[38;2;112;28;6m.\033[38;2;148;78;44m--\033[38;2;138;75;37m-\033[38;2;155;84;50m-\033[38;2;160;93;61m=\033[38;2;172;99;74m=\033[38;2;168;98;73m=\033[38;2;172;97;75m=\033[38;2;173;98;73m=\033[38;2;164;92;67m==\033[38;2;158;81;44m-\033[38;2;163;80;40m-\033[38;2;174;98;63m=\033[38;2;179;97;68m=\033[38;2;180;104;77m=\033[38;2;179;102;72m=\033[38;2;166;84;47m=\033[38;2;171;87;51m=\033[38;2;197;129;98m+\033[38;2;204;131;108m+\033[38;2;178;86;68m=\033[38;2;210;135;122m*\033[38;2;224;165;151m*\033[38;2;221;141;135m*\033[38;2;198;107;81m++\033[38;2;188;105;97m=\033[38;2;153;75;62m-\033[38;2;168;94;81m=\033[38;2;174;98;93m=\033[38;2;130;47;44m:\033[38;2;97;6;8m.\033[38;2;78;1;4m \033[38;2;60;0;0m \033[38;2;67;7;6m \033[38;2;75;13;19m.\033[38;2;59;1;4m .\033[38;2;184;133;115m+\033[38;2;102;19;3m.\033[38;2;118;43;1m:\033[38;2;110;57;22m:\033[38;2;64;4;0m \033[38;2;66;17;6m.\033[38;2;67;26;14m.\033[38;2;47;9;6m \033[38;2;32;1;2m   \033[38;2;34;4;0m \033[38;2;45;29;17m.\033[38;2;77;55;41m:\033[38;2;187;161;160m*\033[38;2;252;251;248m@@@@\033[38;2;253;244;244m@\033[38;2;255;241;242m@@\033[38;2;253;233;236m@@\033[38;2;252;210;209m&\033[38;2;248;211;202m&\033[38;2;252;208;193m&\033[38;2;246;182;160m#\033[38;2;230;165;137m*\033[38;2;227;160;132m*\033[38;2;237;171;145m#\033[38;2;233;166;139m#\033[38;2;242;174;152m#\033[38;2;238;177;149m#\033[38;2;241;179;154m#\033[38;2;251;194;167m&\033[38;2;247;188;157m#\033[38;2;248;200;178m&\033[38;2;214;147;112m*\033[38;2;229;164;133m*\033[38;2;233;180;148m#\033[38;2;255;206;180m&&&\033[38;2;249;205;188m&\033[0m");
        $display("\033[38;2;1;2;4m \033[38;2;98;72;67m-\033[38;2;112;48;37m:\033[38;2;115;42;23m:\033[38;2;106;25;10m.\033[38;2;85;5;0m.\033[38;2;137;86;47m-\033[38;2;129;90;52m-\033[38;2;132;99;46m-\033[38;2;103;36;3m::\033[38;2;100;43;0m:\033[38;2;121;68;3m:\033[38;2;116;52;8m:\033[38;2;185;143;110m+\033[38;2;228;199;165m#\033[38;2;193;151;115m*\033[38;2;149;105;53m=\033[38;2;76;17;1m.\033[38;2;63;1;3m \033[38;2;74;10;6m.\033[38;2;133;84;38m-\033[38;2;116;65;2m:\033[38;2;156;99;44m=\033[38;2;150;96;38m=\033[38;2;208;168;134m*\033[38;2;191;152;111m*\033[38;2;65;17;6m.\033[38;2;66;13;2m.\033[38;2;144;90;66m-\033[38;2;153;89;57m=\033[38;2;249;216;184m&\033[38;2;79;14;12m.\033[38;2;109;34;24m:\033[38;2;124;56;45m:\033[38;2;136;69;43m-\033[38;2;156;99;73m=\033[38;2;153;86;38m--\033[38;2;178;112;76m=\033[38;2;172;99;69m==\033[38;2;158;76;46m-\033[38;2;170;88;57m=\033[38;2;164;89;60m=\033[38;2;160;85;51m=\033[38;2;155;80;42m-\033[38;2;162;82;50m-\033[38;2;152;70;18m-\033[38;2;169;99;72m=\033[38;2;170;98;65m=\033[38;2;168;100;69m=\033[38;2;158;77;28m-\033[38;2;184;108;77m=\033[38;2;181;111;86m=\033[38;2;189;122;96m+\033[38;2;200;111;101m+\033[38;2;163;78;56m-\033[38;2;151;49;34m-\033[38;2;147;70;55m-\033[38;2;110;16;12m.\033[38;2;71;2;3m \033[38;2;52;0;0m \033[38;2;90;46;40m:\033[38;2;129;90;87m-\033[38;2;206;169;170m*\033[38;2;137;112;107m=\033[38;2;85;41;40m:\033[38;2;60;9;8m \033[38;2;45;1;0m  \033[38;2;60;18;17m.\033[38;2;61;2;2m  \033[38;2;204;154;141m*\033[38;2;131;60;32m-\033[38;2;122;61;31m:\033[38;2;98;49;14m:\033[38;2;64;1;0m \033[38;2;82;23;12m.\033[38;2;62;2;0m \033[38;2;91;48;33m:\033[38;2;68;26;8m.\033[38;2;79;53;35m:\033[38;2;69;33;25m.\033[38;2;98;55;48m:\033[38;2;235;220;210m&\033[38;2;254;251;252m@@@\033[38;2;253;241;248m@\033[38;2;255;238;243m@@@@\033[38;2;253;240;247m@@\033[38;2;254;235;241m@@\033[38;2;252;226;214m&\033[38;2;255;198;186m&\033[38;2;245;183;162m#\033[38;2;232;165;137m#\033[38;2;220;154;120m*\033[38;2;224;151;116m*\033[38;2;205;136;95m+\033[38;2;217;148;117m*\033[38;2;236;172;142m#\033[38;2;246;183;154m#\033[38;2;251;196;165m&\033[38;2;254;199;176m&\033[38;2;247;187;160m#\033[38;2;230;164;132m*\033[38;2;224;159;128m*\033[38;2;242;185;156m#\033[38;2;254;200;176m&&\033[38;2;255;204;183m&\033[38;2;250;218;198m&\033[0m");
        $display("\033[38;2;4;4;6m \033[38;2;77;48;44m:\033[38;2;118;56;46m:\033[38;2;109;37;29m:\033[38;2;113;52;32m:\033[38;2;101;30;5m.\033[38;2;104;49;9m:\033[38;2;123;77;21m-\033[38;2;190;156;120m*\033[38;2;157;117;63m=\033[38;2;134;79;11m-\033[38;2;138;92;38m-\033[38;2;120;58;6m:\033[38;2;158;116;67m=\033[38;2;239;209;194m&\033[38;2;250;243;225m@\033[38;2;223;199;169m#\033[38;2;183;148;110m+\033[38;2;89;30;9m.\033[38;2;64;4;3m \033[38;2;67;3;4m \033[38;2;112;54;16m:\033[38;2;137;89;35m-\033[38;2;135;75;11m-\033[38;2;193;162;113m*\033[38;2;221;190;155m#\033[38;2;217;180;148m#\033[38;2;61;8;4m \033[38;2;55;10;5m \033[38;2;64;16;13m.\033[38;2;204;162;139m*\033[38;2;130;91;46m-\033[38;2;207;181;168m#\033[38;2;67;41;20m.\033[38;2;59;12;7m  \033[38;2;145;88;55m-\033[38;2;159;83;58m-\033[38;2;120;36;2m:\033[38;2;158;78;38m--\033[38;2;175;108;79m==\033[38;2;169;98;65m=\033[38;2;179;108;83m=\033[38;2;157;82;39m-\033[38;2;156;78;38m-\033[38;2;159;84;56m-\033[38;2;140;57;7m:\033[38;2;155;80;38m-\033[38;2;161;82;47m-\033[38;2;163;93;55m=\033[38;2;148;61;13m-\033[38;2;195;130;105m+\033[38;2;173;111;78m=\033[38;2;133;48;20m:\033[38;2;125;14;10m.\033[38;2;116;27;20m:\033[38;2;110;44;47m:\033[38;2;78;29;33m.\033[38;2;36;4;2m \033[38;2;27;1;3m \033[38;2;6;2;0m   \033[38;2;2;0;1m  \033[38;2;38;4;6m \033[38;2;70;30;30m.\033[38;2;39;0;0m \033[38;2;45;1;1m \033[38;2;49;5;5m .\033[38;2;129;43;31m:\033[38;2;199;157;138m*\033[38;2;153;98;69m=\033[38;2;119;73;37m-\033[38;2;57;0;0m \033[38;2;64;3;8m \033[38;2;72;30;14m.\033[38;2;77;10;3m.\033[38;2;99;42;2m:\033[38;2;174;137;111m+\033[38;2;236;220;196m&\033[38;2;249;247;239m@\033[38;2;250;253;254m@\033[38;2;255;252;255m@\033[38;2;253;235;240m@\033[38;2;248;221;220m&\033[38;2;254;227;226m@\033[38;2;240;208;203m&\033[38;2;250;216;212m&\033[38;2;252;224;219m&\033[38;2;253;221;223m&@@\033[38;2;249;249;247m@\033[38;2;254;250;252m@\033[38;2;251;229;224m@\033[38;2;247;198;184m&&\033[38;2;255;206;192m&\033[38;2;254;199;177m&\033[38;2;251;194;167m&\033[38;2;218;152;117m*\033[38;2;184;118;69m+\033[38;2;229;162;127m*\033[38;2;235;175;142m#\033[38;2;250;192;164m#\033[38;2;249;195;165m&\033[38;2;255;208;182m&\033[38;2;249;202;175m&\033[38;2;243;182;151m#\033[38;2;221;161;128m*\033[38;2;233;171;140m#\033[38;2;253;202;174m&\033[38;2;254;224;198m&&\033[38;2;253;237;219m@\033[0m");
        $display("\033[38;2;0;4;3m \033[38;2;26;1;0m \033[38;2;64;7;5m \033[38;2;84;11;1m..\033[38;2;86;7;9m.\033[38;2;93;30;7m.\033[38;2;92;15;0m.\033[38;2;142;101;47m=\033[38;2;215;184;158m#\033[38;2;177;144;111m+\033[38;2;157;115;74m=\033[38;2;121;53;3m:\033[38;2;218;191;172m#\033[38;2;254;253;249m@\033[38;2;253;255;243m@\033[38;2;252;234;213m@\033[38;2;188;154;126m*\033[38;2;60;23;7m.\033[38;2;65;8;3m \033[38;2;61;2;4m \033[38;2;75;14;2m.\033[38;2;124;74;31m-\033[38;2;141;80;27m-\033[38;2;166;130;70m+\033[38;2;213;175;136m#\033[38;2;210;176;147m#\033[38;2;84;33;18m.\033[38;2;51;13;6m \033[38;2;45;15;2m \033[38;2;48;1;7m \033[38;2;131;87;71m-\033[38;2;194;159;127m*\033[38;2;234;215;194m&\033[38;2;92;72;57m:\033[38;2;56;3;0m \033[38;2;110;43;33m:\033[38;2;118;54;12m:\033[38;2;148;75;39m-\033[38;2;152;77;37m-\033[38;2;154;81;45m-\033[38;2;171;105;72m=\033[38;2;161;87;51m==\033[38;2;188;112;89m+\033[38;2;170;93;55m==\033[38;2;156;83;50m-\033[38;2;157;79;43m-\033[38;2;162;87;49m=\033[38;2;160;92;58m=\033[38;2;173;109;75m=\033[38;2;153;82;27m-\033[38;2;198;137;109m+\033[38;2;160;92;76m=\033[38;2;75;0;0m \033[38;2;81;12;11m.\033[38;2;64;21;9m.\033[38;2;40;1;2m \033[38;2;2;3;1m \033[38;2;3;2;6m \033[38;2;21;4;2m  \033[38;2;42;3;3m \033[38;2;41;2;2m   \033[38;2;49;4;6m \033[38;2;91;49;45m:\033[38;2;88;41;39m:\033[38;2;51;10;6m \033[38;2;53;1;1m \033[38;2;78;0;2m \033[38;2;130;58;45m-\033[38;2;147;95;70m=\033[38;2;152;99;77m=\033[38;2;100;45;15m:\033[38;2;49;0;0m   \033[38;2;107;63;44m:\033[38;2;255;251;249m@@\033[38;2;251;250;246m@\033[38;2;252;252;247m@\033[38;2;254;243;235m@\033[38;2;246;218;201m&\033[38;2;240;198;178m&\033[38;2;255;218;197m&\033[38;2;224;172;156m#\033[38;2;241;189;171m#\033[38;2;224;169;154m#\033[38;2;218;160;144m*\033[38;2;240;188;175m#\033[38;2;247;216;202m&\033[38;2;255;234;225m@\033[38;2;253;221;210m&&\033[38;2;245;189;168m#\033[38;2;253;202;182m&\033[38;2;255;208;188m&\033[38;2;254;209;187m&\033[38;2;250;189;165m#\033[38;2;228;161;132m*\033[38;2;198;132;97m+\033[38;2;191;120;78m+\033[38;2;208;142;102m*\033[38;2;223;163;131m*\033[38;2;246;190;161m#\033[38;2;241;185;152m#\033[38;2;255;207;177m&\033[38;2;254;210;185m&&\033[38;2;247;188;156m#\033[38;2;234;171;143m#\033[38;2;246;182;153m#\033[38;2;254;206;183m&\033[38;2;253;218;196m&\033[38;2;252;231;213m@\033[0m");
        $display("\033[38;2;1;1;0m \033[38;2;31;5;1m \033[38;2;86;36;26m.\033[38;2;81;14;4m.\033[38;2;93;34;10m.\033[38;2;85;25;8m.\033[38;2;72;1;3m \033[38;2;75;0;6m \033[38;2;139;101;65m=\033[38;2;214;187;160m#\033[38;2;168;133;99m+\033[38;2;160;127;97m+\033[38;2;217;195;174m#\033[38;2;252;252;250m@\033[38;2;254;251;245m@@\033[38;2;113;68;52m-\033[38;2;61;2;2m \033[38;2;65;18;0m.\033[38;2;83;47;20m:\033[38;2;55;6;0m \033[38;2;52;0;2m \033[38;2;83;30;6m.\033[38;2;148;107;68m=\033[38;2;166;129;75m+\033[38;2;171;131;79m+\033[38;2;196;163;125m*\033[38;2;122;65;18m:\033[38;2;52;3;0m \033[38;2;42;5;1m \033[38;2;47;9;3m \033[38;2;53;2;0m  \033[38;2;114;64;43m:\033[38;2;249;222;204m&\033[38;2;85;30;17m.\033[38;2;55;0;0m \033[38;2;123;58;33m:\033[38;2;128;56;15m:\033[38;2;142;68;27m-\033[38;2;157;93;57m=\033[38;2;160;87;53m==\033[38;2;187;115;92m+\033[38;2;189;114;93m+\033[38;2;197;126;106m+\033[38;2;176;108;73m=\033[38;2;152;80;27m-\033[38;2;169;83;53m=\033[38;2;154;78;24m-\033[38;2;181;111;83m=\033[38;2;182;117;84m+\033[38;2;192;124;101m+\033[38;2;196;144;125m*\033[38;2;147;66;41m-\033[38;2;74;0;2m \033[38;2;71;36;16m.\033[38;2;55;5;1m \033[38;2;51;1;0m \033[38;2;47;8;1m \033[38;2;72;38;21m.\033[38;2;104;57;51m:\033[38;2;128;80;71m-\033[38;2;138;85;78m-\033[38;2;157;116;105m=\033[38;2;210;172;163m#\033[38;2;121;71;67m-\033[38;2;50;2;1m \033[38;2;69;1;0m \033[38;2;94;37;30m:\033[38;2;59;0;2m \033[38;2;72;1;7m \033[38;2;93;16;11m.\033[38;2;177;120;106m+\033[38;2;155;97;81m==\033[38;2;120;66;33m-\033[38;2;45;0;0m \033[38;2;47;14;9m \033[38;2;155;106;101m=\033[38;2;251;252;249m@@\033[38;2;255;235;229m@@\033[38;2;253;225;218m&\033[38;2;255;209;194m&\033[38;2;251;194;174m&\033[38;2;245;192;169m#\033[38;2;230;183;153m#\033[38;2;242;195;170m#\033[38;2;249;201;188m&&\033[38;2;247;194;190m&\033[38;2;242;193;188m#\033[38;2;239;191;174m#\033[38;2;225;167;145m#*\033[38;2;236;170;153m#\033[38;2;249;184;162m#\033[38;2;243;182;160m##\033[38;2;232;164;136m*\033[38;2;219;153;121m*\033[38;2;231;166;138m#\033[38;2;221;162;129m*\033[38;2;212;147;117m*\033[38;2;186;120;82m+\033[38;2;222;160;129m*\033[38;2;244;183;155m#\033[38;2;241;184;154m#\033[38;2;248;194;163m#\033[38;2;255;219;190m&\033[38;2;254;214;189m&\033[38;2;253;212;185m&\033[38;2;235;170;143m#\033[38;2;228;163;128m*\033[38;2;252;196;170m&\033[38;2;255;210;191m&\033[38;2;254;233;218m@\033[0m");
        $display("\033[38;2;0;2;1m \033[38;2;31;3;2m \033[38;2;33;2;0m \033[38;2;43;3;3m \033[38;2;46;1;6m \033[38;2;53;2;1m  \033[38;2;79;5;0m.\033[38;2;152;114;88m=\033[38;2;226;194;160m#\033[38;2;239;212;182m&\033[38;2;240;232;203m&\033[38;2;255;249;225m@\033[38;2;245;230;195m&\033[38;2;219;201;158m#\033[38;2;199;168;130m*\033[38;2;74;21;7m.\033[38;2;54;18;9m.\033[38;2;95;63;34m:\033[38;2;83;41;24m:\033[38;2;53;2;6m \033[38;2;48;1;3m \033[38;2;58;0;2m \033[38;2;89;45;3m:\033[38;2;140;97;49m=\033[38;2;167;122;80m+\033[38;2;158;121;78m=\033[38;2;133;84;29m-\033[38;2;89;32;8m.\033[38;2;64;11;10m.\033[38;2;41;9;2m \033[38;2;49;11;8m  \033[38;2;84;39;18m.\033[38;2;79;9;8m.\033[38;2;197;146;122m*\033[38;2;200;159;135m*\033[38;2;78;18;14m.\033[38;2;82;12;9m.\033[38;2;114;36;7m:\033[38;2;151;90;66m=\033[38;2;142;77;38m-\033[38;2;147;76;22m-\033[38;2;163;92;61m=\033[38;2;183;117;92m++\033[38;2;182;115;85m+\033[38;2;175;100;72m=\033[38;2;155;78;24m-\033[38;2;181;113;79m=\033[38;2;187;118;96m++\033[38;2;179;113;80m=\033[38;2;140;76;44m-\033[38;2;178;114;97m+\033[38;2;82;1;4m.\033[38;2;116;51;27m:\033[38;2;199;150;137m*\033[38;2;197;151;144m*\033[38;2;167;130;116m+\033[38;2;160;104;95m=\033[38;2;142;99;85m=\033[38;2;149;95;73m=\033[38;2;109;37;12m:\033[38;2;138;83;65m-\033[38;2;176;115;112m+\033[38;2;163;110;84m=\033[38;2;86;7;0m.\033[38;2;174;127;108m+\033[38;2;69;11;3m.\033[38;2;89;37;20m.\033[38;2;73;3;7m \033[38;2;139;49;40m:\033[38;2;168;106;97m=\033[38;2;134;59;39m-\033[38;2;171;123;107m+\033[38;2;92;31;12m.\033[38;2;62;2;3m \033[38;2;119;57;57m:\033[38;2;251;252;243m@\033[38;2;253;235;228m@\033[38;2;255;214;204m&&\033[38;2;253;213;201m&\033[38;2;254;215;203m&\033[38;2;255;208;193m&\033[38;2;235;173;160m#\033[38;2;231;174;155m#\033[38;2;226;180;157m#\033[38;2;247;196;177m&\033[38;2;255;209;195m&&\033[38;2;254;216;204m&\033[38;2;249;207;183m&\033[38;2;232;179;156m#\033[38;2;194;128;98m++\033[38;2;215;146;120m*\033[38;2;218;154;125m**\033[38;2;214;150;117m*\033[38;2;221;157;124m*\033[38;2;237;173;144m#\033[38;2;249;186;155m#\033[38;2;241;182;148m#\033[38;2;235;175;147m#\033[38;2;238;173;145m#\033[38;2;203;140;99m+\033[38;2;238;176;148m##\033[38;2;240;185;156m#\033[38;2;255;224;196m&\033[38;2;250;210;181m&\033[38;2;255;217;191m&\033[38;2;254;208;182m&\033[38;2;218;154;120m*\033[38;2;213;147;117m*\033[38;2;239;178;156m#\033[38;2;253;239;221m@\033[0m");
        $display("\033[38;2;1;1;1m  \033[38;2;34;0;2m \033[38;2;35;4;0m \033[38;2;54;33;17m.\033[38;2;57;18;8m.\033[38;2;160;123;99m+\033[38;2;222;194;179m#\033[38;2;246;244;240m@\033[38;2;253;253;241m@\033[38;2;252;246;227m@\033[38;2;254;239;212m@\033[38;2;239;220;188m&\033[38;2;245;221;181m&\033[38;2;232;205;176m&\033[38;2;163;132;87m+\033[38;2;101;64;9m:\033[38;2;110;78;38m-\033[38;2;94;51;25m:\033[38;2;52;25;8m.\033[38;2;38;2;3m   \033[38;2;105;45;31m:\033[38;2;104;57;23m:\033[38;2;175;138;90m+\033[38;2;116;61;8m::.\033[38;2;79;19;7m.\033[38;2;91;39;9m.\033[38;2;61;6;1m  \033[38;2;53;13;8m \033[38;2;82;25;24m.\033[38;2;86;12;15m.\033[38;2;138;80;47m-\033[38;2;239;200;175m&\033[38;2;120;69;51m-\033[38;2;71;0;1m \033[38;2;94;26;9m.\033[38;2;117;40;17m:\033[38;2;137;66;40m-\033[38;2;141;63;12m-\033[38;2;134;46;5m:\033[38;2;175;100;69m=\033[38;2;184;119;93m++\033[38;2;155;75;30m-\033[38;2;165;94;51m=\033[38;2;201;145;120m*\033[38;2;211;153;123m*\033[38;2;171;106;79m=\033[38;2;173;107;74m=\033[38;2;177;110;84m=\033[38;2;109;6;2m.\033[38;2;76;1;3m \033[38;2;94;25;13m.\033[38;2;150;83;66m-\033[38;2;158;93;78m=\033[38;2;151;91;73m=\033[38;2;155;89;76m=\033[38;2;131;57;44m-\033[38;2;127;51;32m:\033[38;2;165;90;83m=\033[38;2;193;138;129m+\033[38;2;190;134;126m+\033[38;2;210;161;142m*\033[38;2;191;137;106m+\033[38;2;199;157;141m*\033[38;2;226;178;172m#\033[38;2;85;2;2m.\033[38;2;132;48;37m:\033[38;2;206;135;138m*\033[38;2;131;52;40m:\033[38;2;182;117;101m+\033[38;2;78;0;2m \033[38;2;153;92;81m=\033[38;2;254;251;245m@\033[38;2;252;224;212m&&\033[38;2;251;202;192m&\033[38;2;249;193;181m&\033[38;2;243;195;175m#\033[38;2;234;183;164m#\033[38;2;246;189;170m#\033[38;2;223;166;146m*\033[38;2;219;164;143m*\033[38;2;234;190;163m#\033[38;2;224;179;158m#\033[38;2;252;208;191m&\033[38;2;251;205;188m&\033[38;2;238;196;182m#\033[38;2;245;202;178m&\033[38;2;223;180;155m##\033[38;2;213;156;127m*\033[38;2;199;133;101m+\033[38;2;203;135;103m+\033[38;2;212;151;120m*\033[38;2;238;178;150m#\033[38;2;231;172;142m#\033[38;2;243;180;147m#\033[38;2;250;188;157m#\033[38;2;235;180;149m#\033[38;2;253;201;173m&\033[38;2;217;161;126m*\033[38;2;227;166;134m**\033[38;2;246;182;150m#\033[38;2;236;175;144m#\033[38;2;245;188;157m#\033[38;2;254;209;182m&\033[38;2;253;203;180m&\033[38;2;255;216;187m&\033[38;2;248;191;166m#\033[38;2;208;144;112m*\033[38;2;214;149;119m*\033[38;2;250;203;190m&\033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;51;41;36m.\033[38;2;60;36;31m.\033[38;2;131;115;111m=\033[38;2;226;205;199m&\033[38;2;252;239;234m@\033[38;2;255;250;254m@@\033[38;2;252;252;240m@\033[38;2;253;246;225m@\033[38;2;242;219;190m&\033[38;2;236;207;169m&\033[38;2;252;225;202m&\033[38;2;243;224;194m&\033[38;2;169;131;70m+\033[38;2;149;118;64m=\033[38;2;139;108;71m=\033[38;2;137;103;77m=\033[38;2;45;8;0m \033[38;2;47;19;6m.\033[38;2;34;10;3m \033[38;2;38;17;4m \033[38;2;44;1;0m \033[38;2;125;59;43m:\033[38;2;147;103;58m=\033[38;2;139;88;39m-\033[38;2;105;44;3m:\033[38;2;99;34;0m.\033[38;2;86;26;6m.\033[38;2;77;9;1m.\033[38;2;70;3;0m \033[38;2;114;64;43m:\033[38;2;107;69;46m-\033[38;2;68;10;3m. \033[38;2;62;4;4m \033[38;2;105;37;20m:\033[38;2;84;19;21m.\033[38;2;124;48;36m:\033[38;2;182;135;111m+\033[38;2;95;24;17m.\033[38;2;74;1;7m \033[38;2;121;44;26m:\033[38;2;157;89;57m=\033[38;2;130;46;1m:\033[38;2;136;50;5m:\033[38;2;172;101;71m=\033[38;2;182;116;89m+\033[38;2;171;102;71m=\033[38;2;160;77;24m-\033[38;2;159;80;30m-\033[38;2;212;162;131m*\033[38;2;171;108;77m=\033[38;2;128;50;8m:\033[38;2;173;103;82m=\033[38;2;152;77;51m-\033[38;2;124;37;36m:\033[38;2;193;130;118m+\033[38;2;144;69;55m-\033[38;2;192;130;118m+\033[38;2;228;178;178m#\033[38;2;242;195;181m#\033[38;2;237;187;177m#\033[38;2;225;170;158m#\033[38;2;221;163;152m*\033[38;2;230;171;167m#\033[38;2;210;153;141m*\033[38;2;157;75;70m-\033[38;2;93;19;13m.\033[38;2;232;203;187m&\033[38;2;249;225;212m&\033[38;2;104;31;25m:\033[38;2;97;0;0m.\033[38;2;123;2;1m.\033[38;2;150;60;57m-\033[38;2;124;21;15m.\033[38;2;202;152;125m*\033[38;2;252;254;253m@@&\033[38;2;251;200;183m&\033[38;2;245;175;164m#\033[38;2;242;176;158m#\033[38;2;219;162;134m*\033[38;2;218;161;135m*\033[38;2;216;158;136m*\033[38;2;211;151;127m*\033[38;2;214;160;130m*\033[38;2;188;144;107m+\033[38;2;237;192;164m#\033[38;2;213;166;140m*\033[38;2;216;167;148m*\033[38;2;227;180;162m#\033[38;2;207;165;141m*\033[38;2;235;188;166m#\033[38;2;229;183;159m#\033[38;2;196;144;115m*\033[38;2;189;132;102m+\033[38;2;194;135;105m+\033[38;2;208;144;119m*\033[38;2;216;156;128m*\033[38;2;223;158;126m*\033[38;2;225;163;127m*\033[38;2;226;160;126m*\033[38;2;254;195;168m&\033[38;2;242;185;156m#\033[38;2;250;197;165m&\033[38;2;246;191;162m#\033[38;2;230;170;136m#\033[38;2;229;168;140m#\033[38;2;225;164;133m*\033[38;2;240;180;145m#\033[38;2;234;175;141m#\033[38;2;251;198;167m&\033[38;2;254;213;182m&\033[38;2;248;193;176m&\033[38;2;225;162;129m*\033[38;2;194;121;86m+\033[38;2;243;193;173m#\033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;230;224;225m&\033[38;2;149;141;128m+\033[38;2;227;214;204m&\033[38;2;238;230;217m&\033[38;2;251;249;236m@\033[38;2;248;242;231m@\033[38;2;252;255;237m@\033[38;2;235;216;186m&\033[38;2;236;213;176m&\033[38;2;240;221;186m&\033[38;2;254;249;219m@\033[38;2;248;228;196m&\033[38;2;194;164;119m*\033[38;2;141;107;60m=\033[38;2;174;143;103m+\033[38;2;96;58;31m:\033[38;2;64;18;2m.\033[38;2;46;6;1m \033[38;2;44;9;5m \033[38;2;74;26;16m.\033[38;2;105;61;37m:\033[38;2;216;182;153m#\033[38;2;229;202;168m#\033[38;2;164;130;77m+\033[38;2;108;62;10m:\033[38;2;98;53;7m:\033[38;2;71;34;17m.\033[38;2;63;11;2m.\033[38;2;79;31;27m.\033[38;2;50;0;2m \033[38;2;51;1;6m \033[38;2;49;0;0m  \033[38;2;85;14;6m.\033[38;2;97;33;0m.\033[38;2;107;58;21m:\033[38;2;67;16;0m.\033[38;2;71;36;7m.\033[38;2;65;14;10m.\033[38;2;155;104;78m=\033[38;2;177;130;103m+\033[38;2;138;80;59m-\033[38;2;140;66;37m-\033[38;2;135;69;43m-\033[38;2;142;62;31m-\033[38;2;164;98;54m=\033[38;2;179;120;84m+\033[38;2;215;149;122m*\033[38;2;184;117;83m+\033[38;2;153;73;51m-\033[38;2;197;142;107m+\033[38;2;181;113;82m+\033[38;2;180;108;84m=\033[38;2;162;89;56m=\033[38;2;167;106;82m=\033[38;2;160;90;66m=\033[38;2;114;17;15m.\033[38;2;220;159;143m*\033[38;2;224;167;157m#\033[38;2;156;83;69m-\033[38;2;103;0;0m.\033[38;2;97;2;2m.\033[38;2;113;15;11m.\033[38;2;112;26;22m.\033[38;2;76;3;4m \033[38;2;81;1;1m .\033[38;2;153;89;74m=\033[38;2;254;234;222m@\033[38;2;251;246;226m@\033[38;2;86;9;7m.\033[38;2;103;3;1m..\033[38;2;148;35;32m:\033[38;2;229;190;181m#\033[38;2;254;253;249m@\033[38;2;255;235;220m@\033[38;2;252;222;201m&\033[38;2;249;197;167m&\033[38;2;232;173;152m#\033[38;2;243;180;161m#\033[38;2;216;156;128m*\033[38;2;197;142;111m+\033[38;2;193;138;108m+\033[38;2;196;141;109m+\033[38;2;192;137;108m+\033[38;2;190;135;106m+\033[38;2;199;145;121m*\033[38;2;186;136;107m+\033[38;2;178;126;92m+\033[38;2;170;115;76m=\033[38;2;152;97;67m=\033[38;2;149;82;45m-\033[38;2;152;86;56m-\033[38;2;154;98;67m=\033[38;2;123;60;10m:\033[38;2;133;69;32m-\033[38;2;118;48;6m:\033[38;2;126;45;7m:\033[38;2;174;107;57m=\033[38;2;209;148;116m*\033[38;2;229;162;129m*\033[38;2;249;186;158m#\033[38;2;222;163;123m**\033[38;2;238;180;149m#\033[38;2;239;183;155m#\033[38;2;240;180;156m#\033[38;2;235;173;142m#\033[38;2;243;187;161m#\033[38;2;234;166;136m#\033[38;2;244;187;160m#\033[38;2;252;206;178m&\033[38;2;238;184;168m#\033[38;2;246;193;171m#\033[38;2;249;191;180m#\033[38;2;182;102;73m=\033[38;2;157;82;53m-\033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;235;233;233m@\033[38;2;221;216;203m&\033[38;2;245;228;215m&\033[38;2;253;239;222m@@\033[38;2;248;236;217m@\033[38;2;229;206;175m&\033[38;2;241;225;195m&\033[38;2;249;234;206m@\033[38;2;236;206;176m&\033[38;2;199;168;139m*\033[38;2;183;148;113m+\033[38;2;196;163;135m*\033[38;2;119;73;38m-\033[38;2;52;2;0m  \033[38;2;57;1;8m \033[38;2;104;63;18m:\033[38;2;202;163;134m*\033[38;2;244;237;225m@\033[38;2;253;246;227m@\033[38;2;245;226;192m&\033[38;2;167;127;54m+\033[38;2;123;81;18m-\033[38;2;122;70;22m-\033[38;2;77;18;5m.\033[38;2;56;2;0m    \033[38;2;88;20;6m.\033[38;2;113;72;4m:\033[38;2;198;157;123m*\033[38;2;204;164;136m*\033[38;2;184;148;108m+\033[38;2;127;73;3m-\033[38;2;93;22;4m.\033[38;2;77;1;3m \033[38;2;60;0;2m \033[38;2;50;2;0m \033[38;2;111;45;46m:\033[38;2;84;17;3m.\033[38;2;77;1;0m \033[38;2;100;26;16m.\033[38;2;91;1;4m..\033[38;2;88;0;2m.\033[38;2;129;39;22m:\033[38;2;120;22;4m.\033[38;2;106;3;1m.\033[38;2;174;105;67m=\033[38;2;205;154;124m*\033[38;2;156;93;53m=\033[38;2;135;39;1m:\033[38;2;124;28;6m:\033[38;2;156;71;41m-\033[38;2;180;107;93m=\033[38;2;108;10;4m.\033[38;2;253;232;216m@\033[38;2;254;250;244m@\033[38;2;249;241;226m@\033[38;2;255;247;233m@\033[38;2;249;216;207m&\033[38;2;253;247;242m@@\033[38;2;246;213;210m&\033[38;2;254;248;241m@\033[38;2;228;179;163m#\033[38;2;182;118;92m+\033[38;2;88;11;4m.\033[38;2;84;1;7m.\033[38;2;135;35;25m:\033[38;2;235;212;198m&\033[38;2;254;255;249m@\033[38;2;255;241;233m@\033[38;2;253;216;215m&\033[38;2;244;190;164m#\033[38;2;229;165;141m*\033[38;2;218;150;124m*\033[38;2;215;155;130m*\033[38;2;226;167;146m#\033[38;2;203;142;106m*\033[38;2;177;117;77m+\033[38;2;183;114;88m+\033[38;2;173;111;77m=\033[38;2;168;105;72m=\033[38;2;164;101;68m=\033[38;2;163;110;73m=\033[38;2;165;103;71m=\033[38;2;138;79;42m-\033[38;2;139;72;31m-\033[38;2;112;43;2m:\033[38;2;84;18;1m.\033[38;2;70;7;5m. \033[38;2;44;2;4m \033[38;2;41;6;2m   \033[38;2;61;1;1m \033[38;2;134;58;12m:\033[38;2;179;120;80m+\033[38;2;224;161;135m*\033[38;2;211;147;119m*\033[38;2;214;153;122m*\033[38;2;219;154;127m*\033[38;2;214;149;126m*\033[38;2;237;181;158m##\033[38;2;214;152;120m*\033[38;2;230;164;142m*\033[38;2;199;137;95m+\033[38;2;217;145;110m*\033[38;2;218;165;142m*\033[38;2;220;156;145m*\033[38;2;146;70;51m-\033[38;2;98;6;2m.\033[38;2;84;0;0m \033[0m");
        $display("\033[38;2;3;3;5m \033[38;2;242;242;242m@@\033[38;2;250;226;204m&\033[38;2;237;213;189m&\033[38;2;246;221;198m&\033[38;2;209;184;156m#\033[38;2;224;200;168m#\033[38;2;206;185;154m#\033[38;2;221;192;162m#\033[38;2;211;190;151m#\033[38;2;150;124;75m=\033[38;2;155;120;76m=\033[38;2;168;124;94m+\033[38;2;171;117;92m+\033[38;2;218;195;141m#\033[38;2;210;178;144m##\033[38;2;235;219;198m&\033[38;2;248;228;195m&&\033[38;2;197;160;100m*\033[38;2;117;56;0m:\033[38;2;183;153;93m+\033[38;2;197;168;125m*\033[38;2;133;92;14m-\033[38;2;180;131;99m+\033[38;2;167;118;82m=\033[38;2;197;152;106m*\033[38;2;199;163;116m*\033[38;2;229;199;161m#\033[38;2;241;210;179m&&\033[38;2;223;189;156m#\033[38;2;160;121;39m=\033[38;2;126;70;10m-\033[38;2;108;48;4m:\033[38;2;92;29;0m.\033[38;2;100;39;11m:\033[38;2;73;18;13m.\033[38;2;68;9;1m.\033[38;2;98;34;21m:\033[38;2;110;59;37m:\033[38;2;109;41;14m:\033[38;2;82;12;9m.\033[38;2;67;4;3m \033[38;2;94;15;6m.\033[38;2;115;35;23m:\033[38;2;133;63;45m-\033[38;2;134;55;25m:\033[38;2;116;22;5m.\033[38;2;105;16;6m.\033[38;2;228;178;161m#\033[38;2;202;140;120m*\033[38;2;157;87;48m-\033[38;2;124;12;4m.\033[38;2;140;54;41m-\033[38;2;103;1;0m.\033[38;2;138;50;43m:\033[38;2;178;93;90m=\033[38;2;105;18;20m.\033[38;2;165;97;89m=\033[38;2;101;28;10m.\033[38;2;109;26;20m.\033[38;2;124;40;32m:\033[38;2;102;7;7m.\033[38;2;106;12;9m.\033[38;2;118;16;20m.\033[38;2;245;181;179m#\033[38;2;251;217;214m&\033[38;2;207;132;124m+\033[38;2;255;242;236m@@@\033[38;2;253;232;219m@\033[38;2;252;229;216m@\033[38;2;249;198;179m&\033[38;2;235;171;153m#\033[38;2;212;149;121m*\033[38;2;229;167;139m#\033[38;2;222;157;135m*\033[38;2;226;163;132m*\033[38;2;206;137;114m+\033[38;2;172;108;66m=\033[38;2;158;76;30m-\033[38;2;183;114;81m+\033[38;2;200;140;116m+\033[38;2;198;137;110m+\033[38;2;180;116;87m+\033[38;2;156;88;53m=\033[38;2;113;32;0m:\033[38;2;84;12;2m.\033[38;2;75;4;0m \033[38;2;41;0;1m  \033[38;2;32;1;0m \033[38;2;35;0;5m \033[38;2;16;2;1m \033[38;2;5;1;3m \033[38;2;14;0;4m \033[38;2;32;5;0m \033[38;2;57;9;4m \033[38;2;80;12;11m.\033[38;2;122;54;4m:\033[38;2;170;100;68m=\033[38;2;198;136;110m+*\033[38;2;212;143;126m*\033[38;2;227;166;146m#\033[38;2;246;185;158m#\033[38;2;215;153;131m*\033[38;2;175;110;57m=\033[38;2;147;62;27m-\033[38;2;96;18;0m.\033[38;2;76;3;2m  \033[38;2;50;5;6m \033[38;2;55;12;7m \033[38;2;46;5;6m \033[0m");
        $display("\033[38;2;2;2;2m \033[38;2;242;242;241m@\033[38;2;255;249;237m@\033[38;2;243;221;202m&\033[38;2;210;181;153m#\033[38;2;195;165;128m*\033[38;2;158;106;64m==\033[38;2;178;149;120m+\033[38;2;169;152;109m+\033[38;2;146;115;76m=\033[38;2;137;91;64m-\033[38;2;203;180;167m#\033[38;2;247;240;222m@\033[38;2;251;254;247m@@\033[38;2;254;250;244m@@\033[38;2;249;248;237m@\033[38;2;188;148;90m+\033[38;2;174;132;69m+\033[38;2;190;143;100m+\033[38;2;208;176;136m*\033[38;2;190;158;105m*\033[38;2;220;186;147m#\033[38;2;236;208;167m&\033[38;2;238;209;170m&\033[38;2;245;212;179m&\033[38;2;253;225;191m&\033[38;2;254;226;192m&&\033[38;2;240;199;157m#\033[38;2;214;170;121m*\033[38;2;197;153;103m*\033[38;2;164;116;41m==\033[38;2;147;100;45m=\033[38;2;100;43;20m:\033[38;2;85;34;14m.\033[38;2;47;0;1m \033[38;2;60;6;3m \033[38;2;94;41;10m:\033[38;2;103;57;20m:\033[38;2;99;45;4m:\033[38;2;105;46;11m:\033[38;2;108;45;25m:\033[38;2;51;1;1m \033[38;2;46;3;0m  \033[38;2;117;47;34m:\033[38;2;130;51;38m:\033[38;2;102;5;6m.\033[38;2;131;28;15m:\033[38;2;192;140;118m+\033[38;2;215;152;134m*\033[38;2;171;106;81m=\033[38;2;110;13;0m.\033[38;2;131;37;12m:\033[38;2;102;3;1m.\033[38;2;94;0;4m.\033[38;2;107;1;1m.\033[38;2;94;10;3m..\033[38;2;156;51;48m-\033[38;2;139;38;32m:\033[38;2;111;3;1m.\033[38;2;100;1;2m..\033[38;2;120;16;13m.\033[38;2;235;200;183m&\033[38;2;253;244;235m@\033[38;2;254;229;218m@&\033[38;2;255;233;211m@\033[38;2;250;205;188m&\033[38;2;245;185;162m#\033[38;2;235;170;148m##\033[38;2;250;192;172m#\033[38;2;247;190;167m#\033[38;2;227;166;138m*\033[38;2;191;118;83m+\033[38;2;187;115;70m+\033[38;2;178;101;51m=\033[38;2;208;147;120m*\033[38;2;213;158;130m*\033[38;2;210;161;138m*\033[38;2;189;126;97m+\033[38;2;170;113;85m=\033[38;2;154;93;69m=\033[38;2;110;44;22m:\033[38;2;74;1;1m \033[38;2;55;4;2m \033[38;2;35;3;1m \033[38;2;31;0;2m \033[38;2;26;2;6m \033[38;2;2;0;1m \033[38;2;0;2;0m \033[38;2;1;0;5m \033[38;2;2;1;2m \033[38;2;31;2;4m  \033[38;2;49;8;3m \033[38;2;69;10;2m.\033[38;2;93;6;0m.\033[38;2;138;71;28m-\033[38;2;188;135;101m+\033[38;2;203;151;123m*\033[38;2;230;177;153m#\033[38;2;205;148;131m*\033[38;2;194;137;111m+\033[38;2;178;114;89m+\033[38;2;75;4;2m \033[38;2;71;2;0m  \033[38;2;73;17;13m.\033[38;2;58;5;2m \033[38;2;48;9;4m \033[38;2;33;6;2m \033[0m");
        $display("\033[38;2;3;2;2m \033[38;2;234;233;231m&\033[38;2;203;178;170m#\033[38;2;179;148;111m+\033[38;2;250;239;214m@\033[38;2;252;244;228m@\033[38;2;241;232;200m&\033[38;2;191;149;109m*\033[38;2;139;97;30m-\033[38;2;152;118;60m=\033[38;2;175;152;111m+\033[38;2;229;214;200m&\033[38;2;255;255;243m@\033[38;2;254;242;224m@\033[38;2;224;204;182m#\033[38;2;192;163;126m*\033[38;2;162;130;90m+\033[38;2;172;142;96m+\033[38;2;183;145;118m+\033[38;2;157;113;91m=\033[38;2;246;224;200m&\033[38;2;251;231;208m@\033[38;2;226;190;155m#\033[38;2;192;159;124m*\033[38;2;169;124;56m+\033[38;2;180;130;68m+\033[38;2;176;126;65m+\033[38;2;197;144;88m+\033[38;2;218;163;121m*\033[38;2;235;187;150m#\033[38;2;224;180;133m#\033[38;2;226;183;140m#\033[38;2;218;182;133m#\033[38;2;203;166;121m*\033[38;2;201;156;131m*\033[38;2;165;129;76m+\033[38;2;130;85;29m-\033[38;2;97;36;11m.\033[38;2;62;3;2m \033[38;2;49;1;4m \033[38;2;43;0;0m \033[38;2;60;1;3m \033[38;2;62;7;1m \033[38;2;117;71;40m-\033[38;2;99;40;0m:\033[38;2;112;60;18m:\033[38;2;107;67;44m:\033[38;2;59;9;11m \033[38;2;39;24;3m.\033[38;2;58;16;10m.\033[38;2;59;3;1m \033[38;2;113;53;41m:\033[38;2;101;13;4m.\033[38;2;92;4;0m.\033[38;2;201;147;114m*\033[38;2;248;224;209m&\033[38;2;187;134;100m+\033[38;2;186;119;94m+\033[38;2;163;93;63m=\033[38;2;146;59;41m-\033[38;2;126;37;23m:\033[38;2;115;16;10m..\033[38;2;106;8;5m.\033[38;2;138;59;47m-\033[38;2;153;68;58m-\033[38;2;193;133;124m+\033[38;2;252;232;228m@\033[38;2;253;252;247m@\033[38;2;248;230;219m@\033[38;2;247;229;222m@\033[38;2;255;232;219m@\033[38;2;254;222;197m&\033[38;2;250;207;175m&\033[38;2;243;188;161m#\033[38;2;246;184;162m#\033[38;2;244;182;157m#\033[38;2;247;187;161m#\033[38;2;251;193;172m&\033[38;2;226;164;140m*\033[38;2;223;158;126m*\033[38;2;200;133;106m+\033[38;2;217;152;128m*\033[38;2;222;159;134m*\033[38;2;230;174;145m#\033[38;2;219;160;138m*\033[38;2;202;136;112m+\033[38;2;139;45;19m:\033[38;2;150;81;55m-\033[38;2;78;5;3m.\033[38;2;73;11;9m.\033[38;2;44;6;5m  \033[38;2;28;0;4m   \033[38;2;1;1;1m     \033[38;2;38;0;3m  \033[38;2;42;5;0m   \033[38;2;83;16;11m.\033[38;2;142;77;64m-\033[38;2;94;12;0m.\033[38;2;110;40;30m:\033[38;2;94;17;8m.\033[38;2;80;0;1m \033[38;2;78;2;2m \033[38;2;93;34;20m.\033[38;2;80;18;9m.\033[38;2;59;12;4m \033[38;2;46;15;6m \033[38;2;66;35;33m.\033[38;2;14;5;5m \033[0m");
        $display("\033[38;2;4;3;1m \033[38;2;129;118;109m=\033[38;2;72;54;35m:\033[38;2;98;58;47m:\033[38;2;83;34;31m.\033[38;2;168;136;128m+\033[38;2;253;241;227m@\033[38;2;248;249;243m@\033[38;2;255;252;242m@\033[38;2;209;194;178m#\033[38;2;196;173;153m*\033[38;2;144;114;77m=\033[38;2;113;83;66m-\033[38;2;64;42;28m.\033[38;2;69;46;35m:\033[38;2;48;18;12m.\033[38;2;40;4;2m \033[38;2;32;3;0m \033[38;2;33;5;1m \033[38;2;45;20;13m.\033[38;2;53;16;10m.\033[38;2;141;109;90m=\033[38;2;175;142;122m+\033[38;2;143;110;62m=\033[38;2;138;102;34m=\033[38;2;159;111;46m=\033[38;2;169;120;58m=\033[38;2;166;126;60m+\033[38;2;194;155;115m*\033[38;2;188;152;94m*\033[38;2;187;145;90m+++\033[38;2;159;123;78m=\033[38;2;126;87;25m-\033[38;2;100;65;7m:\033[38;2;61;15;1m. \033[38;2;39;0;0m \033[38;2;43;3;1m \033[38;2;36;5;2m  \033[38;2;67;4;0m \033[38;2;69;2;1m \033[38;2;145;98;74m=\033[38;2;129;68;14m-\033[38;2;137;89;42m-\033[38;2;118;76;32m-\033[38;2;76;2;1m  \033[38;2;40;3;2m  \033[38;2;49;12;5m \033[38;2;52;4;0m  \033[38;2;124;51;20m:\033[38;2;173;120;89m+\033[38;2;204;147;133m*\033[38;2;215;157;139m*\033[38;2;195;132;117m+\033[38;2;191;125;113m+\033[38;2;203;142;112m*\033[38;2;210;150;130m*\033[38;2;189;119;98m+\033[38;2;201;150;134m*\033[38;2;238;194;184m#\033[38;2;255;247;244m@@\033[38;2;250;226;212m&\033[38;2;255;238;222m@@\033[38;2;248;203;181m&\033[38;2;249;197;173m&\033[38;2;255;193;172m&\033[38;2;244;188;166m#\033[38;2;254;201;179m&\033[38;2;253;195;175m&\033[38;2;249;189;164m#\033[38;2;238;182;157m#\033[38;2;237;179;155m#\033[38;2;238;176;153m#\033[38;2;229;174;147m#\033[38;2;227;168;143m#\033[38;2;238;175;147m#\033[38;2;215;157;133m*\033[38;2;179;116;85m+\033[38;2;137;89;47m-\033[38;2;84;7;0m. \033[38;2;66;15;15m.\033[38;2;52;18;16m.\033[38;2;30;0;0m          \033[38;2;36;1;3m   \033[38;2;62;19;1m.\033[38;2;64;8;0m   \033[38;2;59;19;3m.\033[38;2;60;9;5m \033[38;2;77;6;4m.\033[38;2;96;36;30m:\033[38;2;73;5;2m \033[38;2;85;23;16m.\033[38;2;58;11;6m \033[38;2;51;12;10m \033[38;2;27;2;2m \033[38;2;20;5;6m \033[38;2;1;1;1m \033[0m");
        $display("\033[38;2;1;1;4m \033[38;2;225;225;225m&\033[38;2;249;247;243m@\033[38;2;213;204;196m#\033[38;2;139;116;103m=\033[38;2;92;74;61m-\033[38;2;54;41;31m.\033[38;2;75;57;51m:\033[38;2;38;18;7m \033[38;2;59;42;27m.\033[38;2;38;17;7m \033[38;2;19;7;3m \033[38;2;4;1;0m  \033[38;2;0;2;3m   \033[38;2;2;0;1m  \033[38;2;16;3;5m \033[38;2;31;17;15m \033[38;2;68;42;33m.\033[38;2;87;68;53m:\033[38;2;76;48;22m:\033[38;2;81;53;14m:\033[38;2;62;26;3m.\033[38;2;94;52;24m:\033[38;2;75;32;2m.\033[38;2;80;29;3m.\033[38;2;105;61;8m:\033[38;2;132;93;48m-\033[38;2;136;102;64m=\033[38;2;113;63;24m:\033[38;2;121;69;30m-\033[38;2;105;58;22m:\033[38;2;95;52;23m:\033[38;2;74;28;19m.\033[38;2;40;0;1m \033[38;2;44;2;4m  \033[38;2;73;40;30m.\033[38;2;50;9;7m \033[38;2;96;48;9m:\033[38;2;102;41;6m:\033[38;2;178;131;99m+\033[38;2;142;93;35m-\033[38;2;193;145;104m+\033[38;2;107;49;9m:\033[38;2;102;48;27m:\033[38;2;94;44;38m:\033[38;2;51;11;10m \033[38;2;43;6;4m \033[38;2;46;5;1m \033[38;2;59;21;10m.\033[38;2;41;2;2m \033[38;2;51;3;1m \033[38;2;59;18;3m.\033[38;2;69;9;1m.\033[38;2;117;53;36m:\033[38;2;192;143;120m+\033[38;2;199;146;125m*\033[38;2;186;125;103m+\033[38;2;146;84;42m-\033[38;2;237;190;175m#\033[38;2;251;247;230m@\033[38;2;253;239;239m@\033[38;2;248;212;205m&\033[38;2;254;218;201m&\033[38;2;251;224;213m&\033[38;2;253;208;197m&\033[38;2;234;176;156m#\033[38;2;243;180;155m#\033[38;2;241;184;160m#\033[38;2;250;196;171m&\033[38;2;255;201;178m&\033[38;2;249;194;173m&\033[38;2;252;201;180m&\033[38;2;254;208;187m&&\033[38;2;255;203;179m&\033[38;2;254;199;175m&\033[38;2;255;203;181m&&\033[38;2;200;144;122m*\033[38;2;169;114;77m=\033[38;2;104;36;1m:\033[38;2;81;23;2m.\033[38;2;54;3;0m \033[38;2;40;11;9m \033[38;2;37;0;1m \033[38;2;24;2;4m \033[38;2;9;1;2m \033[38;2;4;0;5m \033[38;2;0;1;0m      \033[38;2;16;0;1m \033[38;2;34;2;0m  \033[38;2;44;1;2m \033[38;2;40;0;0m \033[38;2;45;7;1m \033[38;2;60;21;4m..\033[38;2;44;3;7m \033[38;2;47;0;0m \033[38;2;67;24;6m.\033[38;2;71;9;5m.\033[38;2;65;2;1m  \033[38;2;67;6;3m \033[38;2;56;12;8m \033[38;2;21;3;2m \033[38;2;7;2;0m   \033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;12;6;3m  \033[38;2;5;0;0m \033[38;2;11;3;1m    \033[38;2;2;0;5m \033[38;2;3;1;4m \033[38;2;1;0;2m         \033[38;2;0;1;0m \033[38;2;9;3;2m \033[38;2;7;2;0m  \033[38;2;17;5;2m  \033[38;2;22;3;0m \033[38;2;53;28;24m.\033[38;2;49;22;8m. \033[38;2;31;1;2m \033[38;2;42;0;6m \033[38;2;45;4;2m \033[38;2;154;119;99m=\033[38;2;109;79;46m-\033[38;2;87;42;18m:\033[38;2;61;16;3m.\033[38;2;76;30;7m.\033[38;2;44;0;0m \033[38;2;57;20;5m.\033[38;2;154;121;107m=\033[38;2;75;44;14m.\033[38;2;55;15;7m.\033[38;2;180;154;124m*\033[38;2;129;84;38m-\033[38;2;179;138;102m+\033[38;2;164;114;60m=\033[38;2;202;168;123m*\033[38;2;128;76;14m-\033[38;2;100;32;6m.\033[38;2;130;89;67m-\033[38;2;49;4;0m \033[38;2;32;12;1m \033[38;2;37;3;2m \033[38;2;44;8;8m   \033[38;2;59;26;11m.\033[38;2;41;7;3m \033[38;2;53;31;8m.\033[38;2;43;4;1m \033[38;2;77;0;2m \033[38;2;210;159;143m*\033[38;2;255;248;245m@\033[38;2;254;254;241m@\033[38;2;246;202;199m&\033[38;2;255;222;220m&\033[38;2;242;210;207m&\033[38;2;255;227;212m@\033[38;2;250;205;190m&\033[38;2;248;186;163m#\033[38;2;236;171;145m#\033[38;2;253;195;171m&\033[38;2;254;198;173m&\033[38;2;255;199;174m&&\033[38;2;251;196;176m&\033[38;2;254;204;181m&&\033[38;2;253;208;186m&&\033[38;2;255;217;197m&\033[38;2;238;184;163m#\033[38;2;220;168;145m*\033[38;2;214;152;135m*\033[38;2;89;12;0m.\033[38;2;92;37;12m.\033[38;2;38;2;1m  \033[38;2;37;3;4m   \033[38;2;2;0;1m        \033[38;2;6;1;0m  \033[38;2;46;0;2m     \033[38;2;67;34;14m.\033[38;2;45;2;2m \033[38;2;41;0;0m \033[38;2;50;10;5m \033[38;2;51;14;13m \033[38;2;40;6;5m \033[38;2;14;0;0m \033[38;2;2;3;4m \033[38;2;1;1;3m \033[38;2;0;0;2m   \033[38;2;1;1;1m \033[0m");
        $display("\033[38;2;0;0;0m             \033[38;2;1;1;1m  \033[38;2;0;0;0m     \033[38;2;8;2;2m  \033[38;2;9;1;0m \033[38;2;10;5;2m  \033[38;2;17;1;1m \033[38;2;57;42;39m.\033[38;2;19;6;1m \033[38;2;27;1;0m    \033[38;2;45;22;12m.\033[38;2;94;41;21m:\033[38;2;208;179;154m#\033[38;2;127;94;56m-\033[38;2;59;2;6m \033[38;2;57;8;1m  \033[38;2;127;88;62m-\033[38;2;95;38;9m:\033[38;2;89;31;6m.\033[38;2;186;150;111m*\033[38;2;112;64;11m:\033[38;2;202;169;135m*\033[38;2;230;207;165m&\033[38;2;216;188;148m#\033[38;2;135;93;25m-\033[38;2;124;84;35m-\033[38;2;111;65;42m:\033[38;2;76;33;19m.\033[38;2;48;1;4m \033[38;2;34;2;3m  \033[38;2;46;7;2m \033[38;2;63;16;8m.\033[38;2;50;0;0m \033[38;2;64;4;3m .\033[38;2;176;127;111m+\033[38;2;255;242;237m@\033[38;2;254;235;231m@@\033[38;2;235;188;178m#\033[38;2;255;229;210m@\033[38;2;254;232;214m@&&\033[38;2;241;179;154m#\033[38;2;246;189;162m#\033[38;2;249;193;166m#\033[38;2;252;196;173m&\033[38;2;254;200;174m&\033[38;2;253;202;175m&\033[38;2;255;204;177m&&&\033[38;2;251;198;178m&\033[38;2;254;201;180m&\033[38;2;255;206;185m&\033[38;2;241;188;170m#\033[38;2;224;176;158m#\033[38;2;201;156;134m*\033[38;2;132;81;62m-\033[38;2;55;2;0m \033[38;2;34;13;7m \033[38;2;20;0;2m \033[38;2;0;1;0m  \033[38;2;2;0;1m          \033[38;2;12;4;2m \033[38;2;39;0;0m  \033[38;2;33;7;7m \033[38;2;17;4;4m \033[38;2;10;0;0m  \033[38;2;2;1;1m      \033[38;2;0;0;0m       \033[0m");
        $display("\033[38;2;0;0;0m     \033[38;2;1;1;1m   \033[38;2;2;2;2m \033[38;2;49;49;49m.\033[38;2;23;23;23m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m     \033[38;2;1;1;1m  \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m  \033[38;2;11;0;0m \033[38;2;20;3;3m \033[38;2;53;35;33m.\033[38;2;24;9;6m \033[38;2;15;1;0m    \033[38;2;47;23;10m.\033[38;2;84;56;35m:\033[38;2;171;149;115m+\033[38;2;177;154;122m*\033[38;2;99;56;16m:\033[38;2;69;2;0m \033[38;2;71;10;6m.\033[38;2;107;61;26m:\033[38;2;112;74;25m-\033[38;2;78;12;0m.\033[38;2;101;46;10m:\033[38;2;198;164;127m*\033[38;2;188;156;112m*\033[38;2;182;149;105m+\033[38;2;157;117;72m=\033[38;2;126;83;37m-\033[38;2;99;50;21m:\033[38;2;113;80;62m-\033[38;2;39;1;1m   \033[38;2;38;8;0m \033[38;2;58;17;8m.\033[38;2;76;5;0m.\033[38;2;216;173;149m#\033[38;2;254;236;220m@\033[38;2;255;233;225m@\033[38;2;253;219;204m&\033[38;2;241;190;179m#\033[38;2;255;213;202m&&\033[38;2;253;220;203m&\033[38;2;249;208;190m&\033[38;2;253;195;176m&\033[38;2;249;197;169m&#\033[38;2;246;190;165m##\033[38;2;252;196;173m&\033[38;2;247;190;170m#\033[38;2;253;198;178m&&\033[38;2;252;196;181m&\033[38;2;250;197;179m&\033[38;2;254;202;181m&\033[38;2;248;196;174m&&\033[38;2;227;176;159m#\033[38;2;210;162;145m*\033[38;2;152;109;85m=\033[38;2;56;10;5m \033[38;2;36;9;4m \033[38;2;4;3;1m    \033[38;2;0;0;0m         \033[38;2;3;1;2m  \033[38;2;7;0;0m  \033[38;2;1;1;1m \033[38;2;0;0;0m                \033[0m");
        $display("\033[38;2;0;0;0m  \033[38;2;7;7;7m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;4;4;4m  \033[38;2;5;5;5m \033[38;2;11;11;11m \033[38;2;1;1;1m \033[38;2;0;0;0m                \033[38;2;1;1;1m \033[38;2;3;4;0m \033[38;2;9;10;5m \033[38;2;7;7;2m \033[38;2;18;15;7m \033[38;2;15;6;4m \033[38;2;14;4;3m \033[38;2;25;0;0m \033[38;2;42;4;4m \033[38;2;72;63;39m:\033[38;2;166;139;115m+\033[38;2;167;150;118m+\033[38;2;132;90;48m-\033[38;2;75;9;2m.\033[38;2;96;39;17m:\033[38;2;75;12;7m.\033[38;2;105;49;6m:\033[38;2;177;139;99m+\033[38;2;117;72;15m-\033[38;2;211;168;134m*\033[38;2;183;142;110m+\033[38;2;148;110;60m=\033[38;2;88;40;5m.:\033[38;2;68;28;12m.\033[38;2;39;3;1m  \033[38;2;47;5;2m \033[38;2;80;18;11m.\033[38;2;227;196;188m#\033[38;2;253;247;235m@\033[38;2;252;236;221m@\033[38;2;253;227;210m&\033[38;2;252;207;189m&\033[38;2;255;214;198m&&\033[38;2;254;212;192m&\033[38;2;249;203;180m&\033[38;2;255;206;181m&\033[38;2;252;194;172m&\033[38;2;247;191;166m#\033[38;2;245;189;164m#\033[38;2;246;190;165m#\033[38;2;247;191;166m#\033[38;2;237;182;157m#\033[38;2;245;189;164m#\033[38;2;234;180;154m#\033[38;2;239;181;157m#\033[38;2;233;175;151m#\033[38;2;229;169;145m#\033[38;2;233;177;152m#\033[38;2;248;192;169m#\033[38;2;232;178;157m#\033[38;2;202;155;124m*\033[38;2;224;180;161m#\033[38;2;178;141;125m+\033[38;2;68;31;11m.\033[38;2;27;13;9m \033[38;2;0;2;1m                                   \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m  \033[38;2;1;1;1m  \033[38;2;2;2;2m \033[38;2;0;0;0m                       \033[38;2;17;3;2m \033[38;2;22;1;0m \033[38;2;20;2;2m \033[38;2;23;1;4m \033[38;2;28;3;1m \033[38;2;51;28;10m.\033[38;2;156;125;99m+\033[38;2;167;143;106m+\033[38;2;126;83;38m-\033[38;2;55;2;0m \033[38;2;73;16;4m.\033[38;2;137;86;56m-\033[38;2;112;69;8m:\033[38;2;126;74;14m-\033[38;2;133;87;37m-\033[38;2;107;62;3m:\033[38;2;72;23;10m.\033[38;2;47;4;6m \033[38;2;65;15;3m.\033[38;2;61;5;8m \033[38;2;48;9;1m \033[38;2;154;100;89m=\033[38;2;227;201;184m#\033[38;2;255;243;228m@\033[38;2;250;241;233m@\033[38;2;255;227;213m@\033[38;2;250;208;194m&\033[38;2;239;190;175m#\033[38;2;253;206;188m&&\033[38;2;252;204;181m&\033[38;2;254;201;177m&&\033[38;2;246;192;164m#\033[38;2;249;193;168m#\033[38;2;252;196;171m&\033[38;2;246;190;165m##\033[38;2;254;196;172m&\033[38;2;245;184;160m#\033[38;2;252;192;168m#\033[38;2;237;183;157m##\033[38;2;242;189;163m#\033[38;2;236;182;156m#\033[38;2;227;176;149m#\033[38;2;230;178;157m#\033[38;2;213;157;135m*\033[38;2;198;156;137m*\033[38;2;174;139;119m+\033[38;2;44;5;0m \033[38;2;32;11;1m \033[38;2;16;2;2m  \033[38;2;0;0;0m                                  \033[0m");
        $display("\033[38;2;0;0;0m    \033[38;2;240;240;240m@\033[38;2;255;255;255m@@@\033[38;2;8;8;8m \033[38;2;0;0;0m    \033[38;2;4;4;4m \033[38;2;255;255;255m@@@@\033[38;2;182;182;182m#\033[38;2;0;0;0m                                                                                                    \033[0m");
        $display("\033[38;2;0;0;0m   \033[38;2;7;7;7m \033[38;2;252;252;252m@\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;17;17;17m \033[38;2;1;1;1m \033[38;2;0;0;0m  \033[38;2;11;11;11m \033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;2;2;2m \033[38;2;0;0;0m                                                                                                    \033[0m");
        $display("\033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;154;154;154m+\033[38;2;255;255;255m@@@@@\033[38;2;252;252;252m@\033[38;2;6;6;6m \033[38;2;0;0;0m  \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;249;249;249m@\033[38;2;0;0;0m   \033[38;2;9;9;9m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@@@\033[38;2;252;252;252m@\033[38;2;253;253;253m@\033[38;2;4;4;4m \033[38;2;0;0;0m    \033[38;2;4;4;4m \033[38;2;92;92;92m-\033[38;2;246;246;246m@\033[38;2;250;250;250m@\033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;250;250;250m@\033[38;2;132;132;132m+\033[38;2;3;3;3m \033[38;2;0;0;0m    \033[38;2;2;2;2m \033[38;2;243;243;243m@\033[38;2;249;249;249m@\033[38;2;255;255;255m@@@@@\033[38;2;247;247;247m@\033[38;2;10;10;10m \033[38;2;0;0;0m    \033[38;2;7;7;7m \033[38;2;4;4;4m \033[38;2;242;242;242m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@\033[38;2;250;250;250m@\033[38;2;254;254;254m@\033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;0;0;0m  \033[38;2;1;1;1m  \033[38;2;129;129;129m=\033[38;2;254;254;254m@\033[38;2;255;255;255m@@@@@\033[38;2;244;244;244m@\033[38;2;106;106;106m=\033[38;2;2;2;2m \033[38;2;0;0;0m    \033[38;2;1;1;1m \033[38;2;241;241;241m@\033[38;2;253;253;253m@@\033[38;2;255;255;255m@@@\033[38;2;251;251;251m@\033[38;2;249;249;249m@\033[38;2;16;16;16m \033[38;2;0;0;0m    \033[38;2;2;2;2m \033[38;2;7;7;7m \033[38;2;249;249;249m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@@@@@\033[38;2;250;250;250m@\033[38;2;2;2;2m \033[0m");
        $display("\033[38;2;1;1;2m \033[38;2;0;0;1m  \033[38;2;250;250;250m@\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;8;8;8m \033[38;2;1;1;1m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;7;7;7m \033[38;2;5;5;5m \033[38;2;2;2;2m \033[38;2;244;244;244m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;250;250;250m@\033[38;2;251;251;251m@\033[38;2;250;250;250m@\033[38;2;251;251;251m@\033[38;2;255;255;255m@@@\033[38;2;138;138;138m+\033[38;2;0;0;0m  \033[38;2;69;69;69m:\033[38;2;255;255;255m@@\033[38;2;251;251;251m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@@@\033[38;2;250;250;250m@\033[38;2;3;3;3m  \033[38;2;11;11;11m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;250;250;250m@\033[38;2;251;251;251m@@\033[38;2;255;255;255m@@@\033[38;2;251;251;251m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;251;251;251m@\033[38;2;253;253;253m@\033[38;2;251;251;251m@\033[38;2;255;255;255m@@\033[38;2;254;254;254m@\033[38;2;88;88;88m-\033[38;2;1;1;1m \033[38;2;14;14;14m \033[38;2;116;116;116m=\033[38;2;252;252;252m@\033[38;2;255;255;255m@@\033[38;2;254;254;254m@@\033[38;2;250;250;250m@\033[38;2;248;248;248m@\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@\033[38;2;249;249;249m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;250;250;250m@\033[38;2;248;248;248m@\033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;6;6;6m \033[38;2;255;255;255m@@@@@\033[38;2;254;254;254m@\033[38;2;255;255;255m@@@@\033[38;2;253;253;253m@\033[0m");
        $display("\033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;37;37;37m.\033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;4;4;4m \033[38;2;250;250;250m@\033[38;2;255;255;255m@@@\033[38;2;215;215;215m&\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;214;214;214m&\033[38;2;1;1;1m \033[38;2;0;0;0m  \033[38;2;146;146;146m+\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@\033[38;2;249;249;249m@\033[38;2;3;3;3m \033[38;2;0;0;0m  \033[38;2;5;5;5m \033[38;2;255;255;255m@@@@\033[38;2;188;188;188m#\033[38;2;2;2;2m \033[38;2;239;239;239m@\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;3;3;3m  \033[38;2;252;252;252m@\033[38;2;255;255;255m@@\033[38;2;249;249;249m@\033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;161;161;161m*\033[38;2;0;0;0m   \033[38;2;190;190;190m#\033[38;2;255;255;255m@@@@\033[38;2;3;3;3m \033[38;2;17;17;17m \033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;6;6;6m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;5;5;5m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@@\033[38;2;143;143;143m+\033[38;2;2;2;2m \033[38;2;233;233;233m&\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;7;7;7m \033[38;2;0;0;0m  \033[38;2;3;3;3m \033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@\033[38;2;254;254;254m@\033[38;2;115;115;115m=\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;6;6;6m \033[38;2;220;220;220m&\033[38;2;255;255;255m@@@\033[0m");
        $display("\033[38;2;0;0;0m  \033[38;2;251;251;251m@\033[38;2;255;255;255m@@\033[38;2;252;252;252m@\033[38;2;229;229;229m&\033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;248;248;248m@\033[38;2;255;255;255m@@@@@@\033[38;2;61;61;61m:\033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;4;4;4m \033[38;2;9;9;9m \033[38;2;0;0;0m \033[38;2;6;6;6m \033[38;2;245;245;245m@\033[38;2;255;255;255m@@@\033[38;2;251;251;251m@\033[38;2;0;0;0m \033[38;2;177;177;177m*\033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;1;1;1m \033[38;2;0;0;0m  \033[38;2;3;3;3m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;61;61;61m:\033[38;2;6;6;6m \033[38;2;251;251;251m@\033[38;2;255;255;255m@@@\033[38;2;89;89;89m-\033[38;2;0;0;0m  \033[38;2;1;1;1m \033[38;2;116;116;116m=\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;1;1;1m \033[38;2;5;5;5m \033[38;2;255;255;255m@@@@\033[38;2;3;3;3m \033[38;2;0;0;0m   \033[38;2;252;252;252m@\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;0;0;0m \033[38;2;232;232;232m&\033[38;2;255;255;255m@@@\033[38;2;248;248;248m@\033[38;2;0;0;0m    \033[38;2;255;255;255m@@@@\033[38;2;28;28;28m.\033[38;2;3;3;3m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;157;157;157m*\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;68;68;68m:\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[38;2;0;0;0m \033[38;2;5;5;5m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;3;3;3m \033[38;2;0;0;0m  \033[38;2;2;2;2m \033[38;2;255;255;255m@@@@\033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;253;253;253m@\033[38;2;255;255;255m@@\033[38;2;254;254;254m@\033[38;2;2;2;2m \033[38;2;0;0;0m  \033[38;2;1;1;1m \033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@@\033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;254;254;254m@\033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;10;10;10m \033[38;2;21;21;21m \033[38;2;248;248;248m@\033[38;2;255;255;255m@@@\033[38;2;253;253;253m@\033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;3;3;3m \033[38;2;252;252;252m@\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;218;218;218m&\033[38;2;4;4;4m \033[38;2;125;125;125m=\033[38;2;254;254;254m@\033[38;2;250;250;250m@\033[38;2;255;255;255m@@\033[38;2;241;241;241m@\033[38;2;0;0;0m  \033[38;2;228;228;228m&\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;47;47;47m.\033[38;2;18;18;18m \033[38;2;250;250;250m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@@\033[38;2;252;252;252m@\033[38;2;9;9;9m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;250;250;250m@\033[38;2;255;255;255m@@@\033[38;2;251;251;251m@\033[38;2;6;6;6m \033[38;2;28;28;28m.\033[38;2;246;246;246m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;9;9;9m \033[38;2;255;255;255m@@@\033[38;2;250;250;250m@\033[38;2;203;203;203m#\033[38;2;8;8;8m \033[38;2;163;163;163m*\033[38;2;244;244;244m@\033[38;2;255;255;255m@@@\033[38;2;229;229;229m&\033[38;2;2;2;2m  \033[38;2;208;208;208m&\033[38;2;251;251;251m@\033[38;2;255;255;255m@@\033[38;2;245;245;245m@\033[38;2;53;53;53m:\033[38;2;6;6;6m \033[38;2;248;248;248m@\033[38;2;255;255;255m@@@@\033[38;2;15;15;15m \033[38;2;0;0;0m  \033[38;2;253;253;253m@\033[38;2;255;255;255m@@\033[38;2;251;251;251m@\033[38;2;246;246;246m@\033[38;2;10;10;10m \033[38;2;38;38;38m.\033[38;2;249;249;249m@\033[38;2;255;255;255m@@@\033[38;2;254;254;254m@\033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;246;246;246m@\033[38;2;255;255;255m@@@\033[38;2;252;252;252m@\033[38;2;2;2;2m \033[38;2;0;0;0m    \033[38;2;245;245;245m@\033[38;2;255;255;255m@@\033[38;2;253;253;253m@\033[38;2;197;197;197m#\033[38;2;2;2;2m \033[38;2;0;0;0m  \033[38;2;6;6;6m \033[38;2;200;200;200m#\033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@@@\033[38;2;254;254;254m@\033[38;2;88;88;88m-\033[38;2;4;4;4m \033[38;2;0;0;0m   \033[38;2;3;3;3m \033[38;2;248;248;248m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@@\033[38;2;252;252;252m@\033[38;2;250;250;250m@\033[38;2;2;2;2m \033[38;2;0;0;0m    \033[38;2;44;44;44m.\033[38;2;253;253;253m@@\033[38;2;255;255;255m@@@@@\033[38;2;247;247;247m@\033[38;2;213;213;213m&\033[38;2;0;0;0m     \033[38;2;216;216;216m&\033[38;2;254;254;254m@@\033[38;2;255;255;255m@@@@\033[38;2;253;253;253m@\033[38;2;248;248;248m@\033[38;2;66;66;66m:\033[38;2;0;0;0m    \033[38;2;4;4;4m \033[38;2;251;251;251m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@@\033[38;2;250;250;250m@@\033[38;2;5;5;5m \033[38;2;0;0;0m   \033[38;2;1;1;1m \033[38;2;31;31;31m.\033[38;2;251;251;251m@\033[38;2;255;255;255m@@@@@@\033[38;2;250;250;250m@\033[38;2;228;228;228m&\033[38;2;2;2;2m \033[38;2;0;0;0m    \033[38;2;242;242;242m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@@@@@\033[38;2;251;251;251m@\033[38;2;252;252;252m@\033[38;2;27;27;27m.\033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;1;1;1m   \033[38;2;6;6;6m \033[38;2;4;4;4m \033[38;2;0;0;0m   \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m  \033[38;2;6;6;6m \033[38;2;2;2;2m \033[38;2;0;0;0m      \033[38;2;2;2;2m \033[38;2;4;4;4m \033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;0;0;0m        \033[38;2;4;4;4m \033[38;2;2;2;2m \033[38;2;4;4;4m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;5;5;5m \033[38;2;3;3;3m \033[38;2;0;0;0m       \033[38;2;3;3;3m \033[38;2;6;6;6m \033[38;2;2;2;2m  \033[38;2;4;4;4m \033[38;2;1;1;1m  \033[38;2;2;2;2m \033[38;2;0;0;0m        \033[38;2;2;2;2m  \033[38;2;3;3;3m  \033[38;2;1;1;1m  \033[38;2;0;0;0m        \033[38;2;2;2;2m \033[38;2;1;1;1m  \033[38;2;2;2;2m \033[38;2;5;5;5m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m        \033[38;2;2;2;2m \033[38;2;3;3;3m \033[38;2;4;4;4m  \033[38;2;1;1;1m  \033[38;2;0;0;0m        \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m  \033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;0;0;0m                                                                                                                      \033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;0;0;0m                                                                                                                     \033[0m");
    end
    endtask

    task you_pass_image;
    begin
        $display("\033[38;2;13;7;9m \033[38;2;11;1;4m \033[38;2;15;1;4m \033[38;2;12;1;1m \033[38;2;9;1;0m \033[38;2;12;0;0m \033[38;2;14;0;0m \033[38;2;14;1;3m \033[38;2;13;1;3m \033[38;2;13;1;3m \033[38;2;13;1;3m \033[38;2;15;0;3m \033[38;2;14;4;5m \033[38;2;13;1;5m \033[38;2;20;5;10m \033[38;2;14;3;7m \033[38;2;5;0;1m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;9;9;9m \033[38;2;39;39;39m.\033[38;2;84;77;80m-\033[38;2;21;11;12m \033[38;2;6;0;0m \033[38;2;5;3;1m \033[38;2;4;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;13;1;5m \033[38;2;16;0;5m \033[38;2;24;3;8m \033[38;2;15;2;3m \033[38;2;9;1;0m \033[38;2;12;0;0m \033[38;2;16;2;2m \033[38;2;20;4;7m \033[38;2;17;1;4m \033[38;2;19;3;6m \033[38;2;13;0;2m \033[38;2;11;1;2m \033[38;2;10;0;1m \033[38;2;12;0;4m \033[38;2;16;0;5m \033[38;2;16;3;7m \033[38;2;9;0;3m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;0;0;1m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;4;4;6m \033[38;2;46;40;42m.\033[38;2;23;13;14m \033[38;2;18;13;13m \033[38;2;10;0;1m \033[38;2;5;3;4m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;18;2;3m \033[38;2;25;4;3m \033[38;2;27;7;9m \033[38;2;28;13;16m \033[38;2;15;1;1m \033[38;2;15;1;1m \033[38;2;18;4;4m \033[38;2;17;1;2m \033[38;2;15;1;1m \033[38;2;13;1;3m \033[38;2;7;1;1m \033[38;2;8;0;1m \033[38;2;10;0;1m \033[38;2;11;0;1m \033[38;2;17;2;5m \033[38;2;17;2;5m \033[38;2;12;0;2m \033[38;2;11;1;2m \033[38;2;3;0;1m \033[38;2;1;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;13;4;5m \033[38;2;138;124;123m=\033[38;2;214;204;199m#\033[38;2;77;65;65m:\033[38;2;35;24;28m.\033[38;2;42;33;34m.\033[38;2;10;6;5m \033[38;2;2;0;1m \033[38;2;4;0;1m \033[38;2;4;0;1m \033[38;2;1;1;1m \033[38;2;1;0;5m \033[38;2;2;2;4m \033[38;2;2;2;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;1;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;3m \033[38;2;0;0;2m \033[38;2;3;0;0m \033[38;2;3;0;0m \033[38;2;3;0;0m \033[38;2;3;0;0m \033[38;2;3;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;2;2;4m \033[38;2;2;2;4m \033[38;2;1;1;3m \033[38;2;2;2;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;20;1;5m \033[38;2;21;2;1m \033[38;2;18;0;0m \033[38;2;16;3;5m \033[38;2;13;1;1m \033[38;2;13;0;0m \033[38;2;14;0;0m \033[38;2;11;0;0m \033[38;2;11;0;1m \033[38;2;12;0;2m \033[38;2;12;0;2m \033[38;2;12;0;2m \033[38;2;20;8;10m \033[38;2;28;13;16m \033[38;2;30;18;22m \033[38;2;27;13;13m \033[38;2;18;6;10m \033[38;2;9;0;3m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;17;11;13m \033[38;2;34;24;23m.\033[38;2;148;135;137m+\033[38;2;233;222;226m&\033[38;2;255;250;247m@\033[38;2;182;175;172m*\033[38;2;54;34;35m.\033[38;2;55;43;45m.\033[38;2;32;24;26m.\033[38;2;12;12;12m \033[38;2;4;1;2m \033[38;2;1;3;2m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;2;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;2;0;3m \033[38;2;9;7;10m \033[38;2;33;28;33m.\033[38;2;54;50;57m:\033[38;2;22;20;23m \033[38;2;85;80;84m-\033[38;2;17;12;16m \033[38;2;3;2;5m \033[38;2;2;2;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;20;1;3m \033[38;2;22;0;3m \033[38;2;21;1;2m \033[38;2;17;0;2m \033[38;2;10;0;0m \033[38;2;12;0;0m \033[38;2;13;1;1m \033[38;2;14;0;2m \033[38;2;14;2;4m \033[38;2;14;2;4m \033[38;2;12;2;3m \033[38;2;9;0;1m \033[38;2;9;1;0m \033[38;2;9;0;0m \033[38;2;13;3;4m \033[38;2;19;3;6m \033[38;2;16;1;4m \033[38;2;9;0;5m \033[38;2;2;0;3m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;2;1;1m \033[38;2;20;5;6m \033[38;2;63;43;43m.\033[38;2;155;135;137m+\033[38;2;188;173;168m*\033[38;2;172;156;149m*\033[38;2;220;208;204m&\033[38;2;242;237;233m@\033[38;2;229;229;225m&\033[38;2;130;118;122m=\033[38;2;45;29;35m.\033[38;2;56;40;45m.\033[38;2;45;36;39m.\033[38;2;21;20;20m \033[38;2;3;1;2m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;1;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;1;0;3m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;1;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;1;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;3;1;1m \033[38;2;2;1;1m \033[38;2;6;4;5m \033[38;2;13;8;12m \033[38;2;26;26;25m.\033[38;2;43;43;43m.\033[38;2;37;30;33m.\033[38;2;119;104;111m=\033[38;2;203;193;202m#\033[38;2;252;245;252m@\033[38;2;232;227;235m&\033[38;2;202;192;200m#\033[38;2;36;22;29m.\033[38;2;17;13;15m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;24;6;6m \033[38;2;43;21;24m.\033[38;2;34;13;23m \033[38;2;28;10;19m \033[38;2;19;0;2m \033[38;2;15;0;0m \033[38;2;16;2;2m \033[38;2;17;2;5m \033[38;2;12;0;2m \033[38;2;9;0;1m \033[38;2;8;0;1m \033[38;2;8;0;1m \033[38;2;12;2;1m \033[38;2;14;0;0m \033[38;2;21;2;9m \033[38;2;25;4;13m \033[38;2;27;10;18m \033[38;2;13;2;5m \033[38;2;6;1;3m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;8;0;0m \033[38;2;25;2;6m \033[38;2;51;15;16m.\033[38;2;171;141;139m+\033[38;2;182;157;153m*\033[38;2;152;123;120m+\033[38;2;180;155;153m*\033[38;2;185;162;162m*\033[38;2;218;198;199m#\033[38;2;254;245;246m@\033[38;2;253;250;249m@\033[38;2;202;183;187m#\033[38;2;106;80;87m-\033[38;2;38;13;19m \033[38;2;52;39;43m.\033[38;2;40;39;40m.\033[38;2;2;1;2m \033[38;2;16;16;16m \033[38;2;6;6;6m \033[38;2;5;5;5m \033[38;2;14;14;14m \033[38;2;9;10;9m \033[38;2;3;4;4m \033[38;2;4;4;4m \033[38;2;5;4;4m \033[38;2;6;4;5m \033[38;2;5;3;4m \033[38;2;15;15;15m \033[38;2;6;6;6m \033[38;2;3;3;3m \033[38;2;6;6;6m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;5;4;6m \033[38;2;20;18;21m \033[38;2;25;23;26m \033[38;2;27;25;28m.\033[38;2;25;23;26m \033[38;2;25;23;28m \033[38;2;16;15;21m \033[38;2;16;15;20m \033[38;2;9;9;11m \033[38;2;3;3;5m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;3m \033[38;2;3;1;4m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;5;5;5m \033[38;2;17;16;14m \033[38;2;32;28;27m.\033[38;2;58;47;50m.\033[38;2;50;32;38m.\033[38;2;58;34;42m.\033[38;2;112;81;90m-\033[38;2;182;164;162m*\033[38;2;255;250;245m@\033[38;2;234;223;221m&\033[38;2;211;199;199m#\033[38;2;167;152;156m*\033[38;2;158;143;146m+\033[38;2;138;121;130m=\033[38;2;25;8;19m \033[38;2;26;22;23m \033[38;2;5;1;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;21;2;4m \033[38;2;30;5;10m \033[38;2;37;12;19m \033[38;2;42;21;32m.\033[38;2;18;4;4m \033[38;2;15;1;1m \033[38;2;15;1;1m \033[38;2;12;2;3m \033[38;2;12;2;3m \033[38;2;17;2;7m \033[38;2;10;1;1m \033[38;2;16;8;4m \033[38;2;16;4;6m \033[38;2;15;0;3m \033[38;2;19;1;6m \033[38;2;24;5;11m \033[38;2;22;2;11m \033[38;2;14;0;6m \033[38;2;18;7;13m \033[38;2;2;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;3;1;2m \033[38;2;4;0;0m \033[38;2;10;6;5m \033[38;2;25;1;3m \033[38;2;91;50;54m:\033[38;2;158;129;125m+\033[38;2;169;144;140m+\033[38;2;187;155;158m*\033[38;2;193;157;159m*\033[38;2;191;159;160m*\033[38;2;180;143;144m+\033[38;2;209;183;184m#\033[38;2;242;230;231m@\033[38;2;253;246;249m@\033[38;2;255;253;255m@\033[38;2;251;253;253m@\033[38;2;238;230;232m&\033[38;2;73;57;64m:\033[38;2;39;19;30m.\033[38;2;127;107;118m=\033[38;2;124;107;117m=\033[38;2;122;105;115m=\033[38;2;109;93;103m-\033[38;2;76;67;72m:\033[38;2;107;102;106m=\033[38;2;165;159;163m*\033[38;2;125;120;124m=\033[38;2;124;119;123m=\033[38;2;142;136;140m+\033[38;2;102;96;100m-\033[38;2;54;41;51m.\033[38;2;26;14;24m \033[38;2;38;28;37m.\033[38;2;49;42;49m.\033[38;2;39;29;37m.\033[38;2;65;55;64m:\033[38;2;151;144;151m+\033[38;2;182;177;181m*\033[38;2;188;183;189m#\033[38;2;159;154;160m*\033[38;2;154;149;155m+\033[38;2;152;150;155m+\033[38;2;151;145;151m+\033[38;2;62;52;60m:\033[38;2;58;52;56m:\033[38;2;51;45;49m.\033[38;2;44;42;43m.\033[38;2;32;30;31m.\033[38;2;32;30;31m.\033[38;2;27;21;23m \033[38;2;19;17;18m \033[38;2;30;30;30m.\033[38;2;40;40;40m.\033[38;2;58;54;53m:\033[38;2;68;50;56m:\033[38;2;57;35;40m.\033[38;2;138;120;122m=\033[38;2;230;222;220m&\033[38;2;253;253;250m@\033[38;2;252;252;250m@\033[38;2;249;237;239m@\033[38;2;212;190;195m#\033[38;2;176;156;155m*\033[38;2;164;140;140m+\033[38;2;169;148;145m+\033[38;2;186;167;169m*\033[38;2;174;162;164m*\033[38;2;142;130;132m+\033[38;2;31;14;20m \033[38;2;17;1;9m \033[38;2;8;2;4m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;22;4;4m \033[38;2;22;0;2m \033[38;2;24;1;8m \033[38;2;30;11;16m \033[38;2;12;0;0m \033[38;2;17;2;2m \033[38;2;22;7;7m \033[38;2;15;1;1m \033[38;2;24;10;10m \033[38;2;24;8;9m \033[38;2;15;2;2m \033[38;2;13;2;1m \033[38;2;14;2;4m \033[38;2;17;1;4m \033[38;2;27;11;17m \033[38;2;26;7;13m \033[38;2;21;2;8m \033[38;2;20;5;12m \033[38;2;43;31;37m.\033[38;2;6;2;4m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;5;4;7m \033[38;2;9;0;3m \033[38;2;29;1;3m \033[38;2;69;44;42m.\033[38;2;167;146;143m+\033[38;2;188;162;161m*\033[38;2;187;151;151m*\033[38;2;184;148;148m*\033[38;2;182;147;145m*\033[38;2;177;148;144m*\033[38;2;172;143;142m+\033[38;2;181;159;156m*\033[38;2;207;185;187m#\033[38;2;225;211;211m&\033[38;2;247;238;239m@\033[38;2;247;244;244m@\033[38;2;254;250;251m@\033[38;2;252;248;249m@\033[38;2;254;250;252m@\033[38;2;254;250;251m@\033[38;2;254;248;248m@\033[38;2;249;248;246m@\033[38;2;253;255;254m@\033[38;2;255;253;254m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;253;253;253m@\033[38;2;250;250;250m@\033[38;2;252;252;252m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;253;251;254m@\033[38;2;255;253;255m@\033[38;2;252;250;251m@\033[38;2;252;251;252m@\033[38;2;253;251;252m@\033[38;2;254;252;253m@\033[38;2;250;248;249m@\033[38;2;252;251;251m@\033[38;2;251;254;253m@\033[38;2;254;252;253m@\033[38;2;255;252;253m@\033[38;2;221;216;217m&\033[38;2;207;199;202m#\033[38;2;222;212;215m&\033[38;2;201;190;196m#\033[38;2;175;164;168m*\033[38;2;176;160;166m*\033[38;2;176;155;156m*\033[38;2;174;157;157m*\033[38;2;248;241;240m@\033[38;2;253;251;253m@\033[38;2;248;246;244m@\033[38;2;243;241;239m@\033[38;2;214;203;203m#\033[38;2;209;189;190m#\033[38;2;170;143;145m+\033[38;2;179;146;147m*\033[38;2;180;144;146m+\033[38;2;170;139;140m+\033[38;2;191;170;167m*\033[38;2;180;158;160m*\033[38;2;195;174;175m*\033[38;2;158;138;140m+\033[38;2;36;8;13m \033[38;2;21;5;6m \033[38;2;5;0;1m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;25;3;6m \033[38;2;31;9;12m \033[38;2;22;0;6m \033[38;2;19;0;5m \033[38;2;15;0;3m \033[38;2;15;0;3m \033[38;2;17;2;5m \033[38;2;13;0;1m \033[38;2;16;1;4m \033[38;2;15;1;1m \033[38;2;8;1;0m \033[38;2;5;0;0m \033[38;2;7;1;1m \033[38;2;14;2;4m \033[38;2;20;4;6m \033[38;2;19;0;3m \033[38;2;13;1;1m \033[38;2;10;0;1m \033[38;2;41;29;33m.\033[38;2;50;40;45m.\033[38;2;3;0;2m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;1m \033[38;2;7;1;3m \033[38;2;6;1;5m \033[38;2;4;2;5m \033[38;2;19;8;7m \033[38;2;48;18;20m.\033[38;2;127;95;96m=\033[38;2;166;146;146m+\033[38;2;177;137;142m+\033[38;2;198;163;161m*\033[38;2;191;158;151m*\033[38;2;201;171;168m*\033[38;2;219;195;192m#\033[38;2;223;202;203m&\033[38;2;234;215;219m&\033[38;2;236;219;220m&\033[38;2;242;224;223m&\033[38;2;243;225;223m&\033[38;2;247;229;227m@\033[38;2;247;229;227m@\033[38;2;249;232;229m@\033[38;2;250;234;231m@\033[38;2;242;228;225m&\033[38;2;244;235;230m@\033[38;2;252;248;247m@\033[38;2;248;238;237m@\033[38;2;247;231;231m@\033[38;2;244;229;232m@\033[38;2;254;239;244m@\033[38;2;249;238;244m@\033[38;2;252;241;247m@\033[38;2;253;244;249m@\033[38;2;254;244;248m@\033[38;2;250;241;243m@\033[38;2;255;247;251m@\033[38;2;248;239;244m@\033[38;2;250;239;247m@\033[38;2;247;238;241m@\033[38;2;244;235;238m@\033[38;2;243;232;236m@\033[38;2;246;237;240m@\033[38;2;246;236;239m@\033[38;2;244;234;234m@\033[38;2;251;241;240m@\033[38;2;242;231;231m@\033[38;2;252;242;243m@\033[38;2;254;252;253m@\033[38;2;255;252;255m@\033[38;2;253;242;241m@\033[38;2;254;240;238m@\033[38;2;255;244;242m@\033[38;2;247;226;225m&\033[38;2;239;215;214m&\033[38;2;214;188;189m#\033[38;2;197;171;170m*\033[38;2;158;133;129m+\033[38;2;171;143;142m+\033[38;2;191;163;163m*\033[38;2;176;148;149m*\033[38;2;199;170;175m*\033[38;2;203;177;182m#\033[38;2;196;177;179m#\033[38;2;164;139;143m+\033[38;2;167;151;153m*\033[38;2;125;105;112m=\033[38;2;60;39;47m.\033[38;2;23;8;15m \033[38;2;6;6;7m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;4;2;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;23;3;5m \033[38;2;20;0;2m \033[38;2;26;3;10m \033[38;2;41;24;28m.\033[38;2;12;2;3m \033[38;2;11;1;2m \033[38;2;12;2;3m \033[38;2;13;1;3m \033[38;2;15;3;5m \033[38;2;21;7;7m \033[38;2;8;3;1m \033[38;2;4;0;0m \033[38;2;8;0;1m \033[38;2;17;2;5m \033[38;2;17;1;2m \033[38;2;20;1;3m \033[38;2;18;4;4m \033[38;2;11;1;2m \033[38;2;15;5;9m \033[38;2;55;49;52m.\033[38;2;10;5;9m \033[38;2;2;2;4m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;3;3;5m \033[38;2;9;1;1m \033[38;2;64;44;44m.\033[38;2;130;101;103m=\033[38;2;187;163;163m*\033[38;2;189;164;160m*\033[38;2;188;164;159m*\033[38;2;167;135;126m+\033[38;2;198;171;164m*\033[38;2;217;189;185m#\033[38;2;240;221;214m&\033[38;2;238;219;215m&\033[38;2;230;210;209m&\033[38;2;238;218;217m&\033[38;2;240;220;221m&\033[38;2;248;228;229m@\033[38;2;252;232;233m@\033[38;2;254;234;235m@\033[38;2;255;235;237m@\033[38;2;253;238;235m@\033[38;2;253;242;235m@\033[38;2;255;249;243m@\033[38;2;249;236;234m@\033[38;2;251;234;234m@\033[38;2;254;235;237m@\033[38;2;254;238;239m@\033[38;2;249;237;237m@\033[38;2;251;239;239m@\033[38;2;252;240;240m@\033[38;2;249;238;242m@\033[38;2;244;234;235m@\033[38;2;247;237;238m@\033[38;2;240;229;233m&\033[38;2;246;234;238m@\033[38;2;246;234;238m@\033[38;2;245;234;238m@\033[38;2;245;234;238m@\033[38;2;238;228;231m&\033[38;2;236;222;227m&\033[38;2;245;229;232m@\033[38;2;240;224;225m&\033[38;2;242;227;228m&\033[38;2;249;229;230m@\033[38;2;229;210;209m&\033[38;2;231;211;210m&\033[38;2;225;205;204m&\033[38;2;204;182;182m#\033[38;2;189;162;159m*\033[38;2;168;138;135m+\033[38;2;159;128;125m+\033[38;2;141;109;106m=\033[38;2;148;116;114m=\033[38;2;175;147;146m+\033[38;2;190;161;163m*\033[38;2;186;160;164m*\033[38;2;187;165;168m*\033[38;2;184;161;164m*\033[38;2;183;162;166m*\033[38;2;204;185;189m#\033[38;2;201;186;188m#\033[38;2;170;151;155m*\033[38;2;26;7;13m \033[38;2;27;18;23m \033[38;2;3;3;5m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;3;1;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[0m");
        $display("\033[38;2;20;1;1m \033[38;2;27;9;9m \033[38;2;22;1;5m \033[38;2;26;9;15m \033[38;2;13;1;3m \033[38;2;10;0;0m \033[38;2;12;4;1m \033[38;2;12;0;2m \033[38;2;14;0;2m \033[38;2;14;2;4m \033[38;2;8;0;1m \033[38;2;6;0;0m \033[38;2;12;2;3m \033[38;2;12;0;2m \033[38;2;16;0;3m \033[38;2;20;3;6m \033[38;2;17;1;2m \033[38;2;10;0;1m \033[38;2;24;13;15m \033[38;2;78;67;73m:\033[38;2;35;33;38m.\033[38;2;7;5;10m \033[38;2;1;1;3m \033[38;2;2;0;3m \033[38;2;2;0;3m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;7;0;0m \033[38;2;10;0;0m \033[38;2;17;0;0m \033[38;2;44;13;11m \033[38;2;93;52;53m:\033[38;2;150;121;117m=\033[38;2;186;160;154m*\033[38;2;214;190;182m#\033[38;2;225;202;194m&\033[38;2;230;205;198m&\033[38;2;225;205;195m&\033[38;2;226;206;196m&\033[38;2;230;209;201m&\033[38;2;233;210;205m&\033[38;2;247;224;218m&\033[38;2;254;232;226m@\033[38;2;252;229;223m@\033[38;2;255;234;228m@\033[38;2;254;240;231m@\033[38;2;252;240;231m@\033[38;2;252;234;224m@\033[38;2;255;238;231m@\033[38;2;248;231;226m@\033[38;2;254;233;230m@\033[38;2;252;236;237m@\033[38;2;245;233;224m@\033[38;2;243;230;224m&\033[38;2;248;235;232m@\033[38;2;234;219;219m&\033[38;2;239;224;227m&\033[38;2;237;220;226m&\033[38;2;237;221;224m&\033[38;2;240;225;227m&\033[38;2;238;222;225m&\033[38;2;236;220;223m&\033[38;2;239;223;226m&\033[38;2;239;223;226m&\033[38;2;239;223;224m&\033[38;2;240;222;222m&\033[38;2;236;218;218m&\033[38;2;238;220;220m&\033[38;2;228;204;204m&\033[38;2;200;176;172m#\033[38;2;197;168;165m*\033[38;2;205;177;168m#\033[38;2;192;163;155m*\033[38;2;184;154;144m*\033[38;2;154;124;114m+\033[38;2;135;102;93m=\033[38;2;134;101;90m=\033[38;2;164;131;124m+\033[38;2;172;138;141m+\033[38;2;189;158;164m*\033[38;2;175;146;150m+\033[38;2;183;160;166m*\033[38;2;217;196;204m#\033[38;2;207;187;196m#\033[38;2;182;165;171m*\033[38;2;131;113;125m=\033[38;2;35;13;28m \033[38;2;25;9;18m \033[38;2;4;4;4m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[0m");
        $display("\033[38;2;41;21;22m.\033[38;2;33;12;16m \033[38;2;22;0;5m \033[38;2;25;6;10m \033[38;2;15;2;2m \033[38;2;19;5;5m \033[38;2;16;3;3m \033[38;2;14;1;4m \033[38;2;20;4;7m \033[38;2;15;0;3m \033[38;2;12;5;5m \033[38;2;6;0;0m \033[38;2;7;0;0m \033[38;2;16;4;6m \033[38;2;25;6;8m \033[38;2;27;4;10m \033[38;2;22;2;3m \033[38;2;24;10;13m \033[38;2;17;1;6m \033[38;2;53;42;50m.\033[38;2;55;49;57m:\033[38;2;3;2;7m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;0;0m \033[38;2;6;0;2m \033[38;2;7;1;1m \033[38;2;32;6;4m \033[38;2;73;29;30m.\033[38;2;191;172;168m*\033[38;2;236;218;208m&\033[38;2;234;216;211m&\033[38;2;231;213;203m&\033[38;2;230;212;200m&\033[38;2;229;207;192m&\033[38;2;227;205;188m&\033[38;2;221;197;186m#\033[38;2;226;201;196m&\033[38;2;237;213;208m&\033[38;2;248;223;218m&\033[38;2;248;223;218m&\033[38;2;251;227;222m@\033[38;2;254;234;226m@\033[38;2;252;232;224m@\033[38;2;253;229;222m@\033[38;2;254;235;226m@\033[38;2;254;236;227m@\033[38;2;252;231;228m@\033[38;2;242;223;219m&\033[38;2;241;222;214m&\033[38;2;240;221;214m&\033[38;2;245;228;221m&\033[38;2;231;211;211m&\033[38;2;235;216;220m&\033[38;2;235;216;222m&\033[38;2;231;212;216m&\033[38;2;230;212;214m&\033[38;2;228;209;211m&\033[38;2;229;210;212m&\033[38;2;233;214;216m&\033[38;2;231;212;214m&\033[38;2;233;215;215m&\033[38;2;225;205;204m&\033[38;2;225;209;206m&\033[38;2;233;212;211m&\033[38;2;228;208;207m&\033[38;2;229;205;201m&\033[38;2;229;206;200m&\033[38;2;217;191;185m#\033[38;2;190;159;154m*\033[38;2;194;165;157m*\033[38;2;180;151;143m*\033[38;2;190;160;154m*\033[38;2;186;159;150m*\033[38;2;171;142;139m+\033[38;2;196;160;167m*\033[38;2;195;162;170m*\033[38;2;176;148;157m*\033[38;2;156;133;141m+\033[38;2;143;125;131m+\033[38;2;169;153;161m*\033[38;2;173;158;168m*\033[38;2;77;59;72m:\033[38;2;22;14;26m \033[38;2;3;2;8m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;4;2;3m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;19;1;1m \033[38;2;21;1;6m \033[38;2;21;0;4m \033[38;2;25;5;8m \033[38;2;19;7;9m \033[38;2;14;2;4m \033[38;2;11;0;1m \033[38;2;10;0;1m \033[38;2;11;1;2m \033[38;2;12;1;3m \033[38;2;12;0;2m \033[38;2;9;0;0m \033[38;2;9;0;1m \033[38;2;11;1;2m \033[38;2;20;5;10m \033[38;2;29;11;13m \033[38;2;22;4;12m \033[38;2;27;6;18m \033[38;2;58;46;55m.\033[38;2;76;68;76m:\033[38;2;78;66;76m:\033[38;2;10;5;11m \033[38;2;4;4;6m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;0;0m \033[38;2;1;1;0m \033[38;2;15;0;3m \033[38;2;36;0;1m \033[38;2;129;106;100m=\033[38;2;239;207;211m&\033[38;2;234;215;204m&\033[38;2;233;209;204m&\033[38;2;229;208;199m&\033[38;2;225;203;192m&\033[38;2;230;209;202m&\033[38;2;231;208;198m&\033[38;2;223;198;182m#\033[38;2;223;195;181m#\033[38;2;239;212;197m&\033[38;2;250;219;204m&\033[38;2;251;219;204m&\033[38;2;254;223;208m&\033[38;2;253;229;211m@\033[38;2;252;229;214m@\033[38;2;254;228;217m@\033[38;2;254;230;218m@\033[38;2;241;218;206m&\033[38;2;245;223;211m&\033[38;2;250;229;217m@\033[38;2;241;223;208m&\033[38;2;248;229;219m@\033[38;2;240;222;216m&\033[38;2;229;212;206m&\033[38;2;234;219;213m&\033[38;2;236;220;221m&\033[38;2;236;220;220m&\033[38;2;236;221;219m&\033[38;2;234;219;222m&\033[38;2;235;221;222m&\033[38;2;230;215;217m&\033[38;2;226;212;212m&\033[38;2;230;215;214m&\033[38;2;228;212;212m&\033[38;2;221;207;207m&\033[38;2;219;201;200m#\033[38;2;228;208;207m&\033[38;2;220;196;192m#\033[38;2;200;177;171m#\033[38;2;224;201;194m#\033[38;2;199;175;169m*\033[38;2;205;179;172m#\033[38;2;188;160;154m*\033[38;2;181;153;148m*\033[38;2;171;140;136m+\033[38;2;166;137;133m+\033[38;2;164;141;138m+\033[38;2;153;126;128m+\033[38;2;148;126;130m+\033[38;2;206;190;193m#\033[38;2;218;201;204m#\033[38;2;98;72;78m-\033[38;2;21;5;10m \033[38;2;17;7;11m \033[38;2;6;3;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;5;1;2m \033[38;2;6;2;3m \033[38;2;6;2;3m \033[38;2;3;0;1m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;24;4;5m \033[38;2;22;1;6m \033[38;2;32;10;15m \033[38;2;42;22;24m.\033[38;2;13;3;4m \033[38;2;11;1;2m \033[38;2;11;1;2m \033[38;2;11;1;2m \033[38;2;12;2;3m \033[38;2;13;1;3m \033[38;2;13;3;4m \033[38;2;10;0;1m \033[38;2;12;2;3m \033[38;2;14;1;3m \033[38;2;21;5;11m \033[38;2;16;4;4m \033[38;2;11;0;3m \033[38;2;12;1;9m \033[38;2;21;8;17m \033[38;2;32;20;29m \033[38;2;67;57;66m:\033[38;2;26;21;27m \033[38;2;3;2;7m \033[38;2;0;0;3m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;3;1;4m \033[38;2;10;5;3m \033[38;2;28;0;1m \033[38;2;111;80;77m-\033[38;2;208;189;182m#\033[38;2;253;234;232m@\033[38;2;232;213;202m&\033[38;2;233;206;199m&\033[38;2;221;196;189m#\033[38;2;216;196;189m#\033[38;2;229;203;197m&\033[38;2;221;190;187m#\033[38;2;233;202;192m&\033[38;2;224;196;181m#\033[38;2;237;209;195m&\033[38;2;240;211;195m&\033[38;2;243;211;196m&\033[38;2;250;217;203m&\033[38;2;252;221;205m&\033[38;2;250;222;208m&\033[38;2;245;218;201m&\033[38;2;243;216;199m&\033[38;2;253;226;209m&\033[38;2;238;212;196m&\033[38;2;227;201;185m#\033[38;2;225;202;184m#\033[38;2;221;197;185m#\033[38;2;208;183;177m#\033[38;2;216;195;188m#\033[38;2;220;202;195m#\033[38;2;223;205;205m&\033[38;2;222;207;202m&\033[38;2;211;198;192m#\033[38;2;214;198;199m#\033[38;2;232;216;219m&\033[38;2;227;211;213m&\033[38;2;230;216;214m&\033[38;2;235;222;215m&\033[38;2;232;217;217m&\033[38;2;221;207;207m&\033[38;2;214;196;192m#\033[38;2;208;188;187m#\033[38;2;212;188;184m#\033[38;2;210;186;182m#\033[38;2;202;178;174m#\033[38;2;188;164;159m*\033[38;2;199;176;170m#\033[38;2;208;186;180m#\033[38;2;190;169;164m*\033[38;2;181;156;152m*\033[38;2;187;163;159m*\033[38;2;179;160;156m*\033[38;2;181;156;158m*\033[38;2;167;147;150m+\033[38;2;227;217;218m&\033[38;2;213;198;201m#\033[38;2;45;24;29m.\033[38;2;30;25;26m.\033[38;2;4;0;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;4;0;1m \033[38;2;6;0;2m \033[38;2;14;8;10m \033[38;2;19;15;16m \033[38;2;3;1;2m \033[0m");
        $display("\033[38;2;30;10;11m \033[38;2;21;1;5m \033[38;2;20;1;2m \033[38;2;23;4;6m \033[38;2;12;0;2m \033[38;2;8;0;0m \033[38;2;5;1;0m \033[38;2;7;1;1m \033[38;2;10;0;1m \033[38;2;11;1;2m \033[38;2;10;1;1m \033[38;2;10;0;1m \033[38;2;13;1;3m \033[38;2;16;1;4m \033[38;2;18;2;5m \033[38;2;17;2;5m \033[38;2;12;0;2m \033[38;2;14;3;11m \033[38;2;20;3;19m \033[38;2;38;24;37m.\033[38;2;94;87;95m-\033[38;2;63;63;65m:\033[38;2;9;4;10m \033[38;2;3;3;5m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;5;1;2m \033[38;2;24;16;14m \033[38;2;37;6;4m \033[38;2;183;167;160m*\033[38;2;240;220;214m&\033[38;2;211;191;183m#\033[38;2;181;153;141m*\033[38;2;109;65;58m:\033[38;2;102;63;56m:\033[38;2;164;136;128m+\033[38;2;219;196;183m#\033[38;2;248;229;220m@\033[38;2;240;219;210m&\033[38;2;251;225;214m&\033[38;2;235;207;195m&\033[38;2;240;213;198m&\033[38;2;241;209;194m&\033[38;2;250;218;203m&\033[38;2;253;220;205m&\033[38;2;251;222;206m&\033[38;2;240;212;195m&\033[38;2;231;205;188m&\033[38;2;230;204;187m&\033[38;2;225;200;181m#\033[38;2;221;196;176m#\033[38;2;216;191;171m#\033[38;2;223;198;183m#\033[38;2;232;205;197m&\033[38;2;238;219;210m&\033[38;2;232;213;209m&\033[38;2;233;216;212m&\033[38;2;236;221;216m&\033[38;2;238;227;215m&\033[38;2;250;238;238m@\033[38;2;246;232;232m@\033[38;2;232;216;217m&\033[38;2;236;223;217m&\033[38;2;238;228;219m&\033[38;2;237;223;220m&\033[38;2;238;224;223m&\033[38;2;242;224;222m&\033[38;2;231;211;210m&\033[38;2;210;187;184m#\033[38;2;209;185;181m#\033[38;2;211;187;185m#\033[38;2;210;186;186m#\033[38;2;206;182;180m#\033[38;2;201;177;176m#\033[38;2;210;186;189m#\033[38;2;201;177;175m#\033[38;2;168;145;139m+\033[38;2;131;108;103m=\033[38;2;153;139;134m+\033[38;2;201;192;189m#\033[38;2;226;212;212m&\033[38;2;89;76;80m-\033[38;2;34;24;28m.\033[38;2;6;6;8m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;2m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;0;1m \033[38;2;11;2;3m \033[38;2;25;16;17m \033[38;2;13;4;5m \033[38;2;5;1;2m \033[38;2;3;1;2m \033[0m");
        $display("\033[38;2;18;4;4m \033[38;2;19;1;3m \033[38;2;12;0;2m \033[38;2;17;3;3m \033[38;2;10;0;1m \033[38;2;10;0;1m \033[38;2;10;0;1m \033[38;2;11;0;1m \033[38;2;11;0;4m \033[38;2;11;0;4m \033[38;2;9;0;3m \033[38;2;12;1;5m \033[38;2;17;4;11m \033[38;2;22;7;14m \033[38;2;19;4;9m \033[38;2;12;1;5m \033[38;2;6;0;2m \033[38;2;8;0;11m \033[38;2;26;11;30m \033[38;2;22;6;25m \033[38;2;35;22;39m.\033[38;2;85;78;94m-\033[38;2;19;15;30m \033[38;2;4;3;6m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;14;10;10m \033[38;2;48;31;29m.\033[38;2;122;99;93m=\033[38;2;227;223;211m&\033[38;2;238;220;210m&\033[38;2;244;226;215m&\033[38;2;235;216;201m&\033[38;2;146;101;92m=\033[38;2;70;37;35m.\033[38;2;66;54;55m:\033[38;2;61;50;55m:\033[38;2;69;45;43m:\033[38;2;86;41;37m:\033[38;2;234;208;198m&\033[38;2;255;238;228m@\033[38;2;242;214;202m&\033[38;2;237;211;194m&\033[38;2;242;216;198m&\033[38;2;252;214;201m&\033[38;2;243;220;202m&\033[38;2;249;213;202m&\033[38;2;247;216;204m&\033[38;2;251;221;210m&\033[38;2;255;235;224m@\033[38;2;241;213;202m&\033[38;2;214;192;170m#\033[38;2;168;136;125m+\033[38;2;134;98;92m=\033[38;2;148;115;109m=\033[38;2;153;123;121m+\033[38;2;45;16;17m \033[38;2;80;54;55m:\033[38;2;50;24;25m.\033[38;2;94;59;55m:\033[38;2;130;101;97m=\033[38;2;203;191;183m#\033[38;2;237;224;215m&\033[38;2;241;217;210m&\033[38;2;245;227;223m&\033[38;2;244;226;224m&\033[38;2;247;229;229m@\033[38;2;253;235;235m@\033[38;2;249;231;231m@\033[38;2;245;226;232m&\033[38;2;246;227;229m&\033[38;2;240;222;222m&\033[38;2;239;221;221m&\033[38;2;240;222;222m&\033[38;2;245;227;227m&\033[38;2;240;222;222m&\033[38;2;224;206;206m&\033[38;2;182;166;166m*\033[38;2;231;217;217m&\033[38;2;252;245;246m@\033[38;2;115;99;105m=\033[38;2;66;57;60m:\033[38;2;22;20;21m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;7;3;4m \033[38;2;15;5;6m \033[38;2;32;20;22m \033[38;2;22;7;10m \033[38;2;6;2;3m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;38;18;20m \033[38;2;36;7;12m \033[38;2;21;0;5m \033[38;2;23;4;6m \033[38;2;15;0;3m \033[38;2;15;0;3m \033[38;2;15;0;3m \033[38;2;12;0;2m \033[38;2;12;1;5m \033[38;2;13;2;6m \033[38;2;8;1;3m \033[38;2;11;0;4m \033[38;2;16;3;10m \033[38;2;20;5;12m \033[38;2;21;6;11m \033[38;2;20;8;12m \033[38;2;13;1;5m \033[38;2;28;14;27m \033[38;2;48;29;49m.\033[38;2;40;24;43m.\033[38;2;34;23;40m.\033[38;2;78;72;84m:\033[38;2;34;30;45m.\033[38;2;5;4;7m \033[38;2;2;1;6m \033[38;2;1;1;1m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;14;3;2m \033[38;2;75;51;49m:\033[38;2;215;199;190m#\033[38;2;237;224;213m&\033[38;2;238;211;203m&\033[38;2;250;232;218m@\033[38;2;253;234;225m@\033[38;2;254;249;240m@\033[38;2;232;209;194m&\033[38;2;130;103;92m=\033[38;2;51;25;14m.\033[38;2;49;15;11m \033[38;2;109;75;65m-\033[38;2;240;216;209m&\033[38;2;251;224;217m&\033[38;2;228;198;187m#\033[38;2;223;190;175m#\033[38;2;227;197;181m#\033[38;2;236;200;186m&\033[38;2;235;206;192m&\033[38;2;235;211;197m&\033[38;2;247;223;209m&\033[38;2;239;203;194m&\033[38;2;164;112;101m=\033[38;2;72;7;6m.\033[38;2;73;46;46m:\033[38;2;61;45;50m.\033[38;2;46;37;42m.\033[38;2;48;46;41m.\033[38;2;52;42;40m.\033[38;2;75;51;55m:\033[38;2;72;37;43m.\033[38;2;183;158;157m*\033[38;2;237;230;218m&\033[38;2;252;242;232m@\033[38;2;250;233;226m@\033[38;2;241;223;216m&\033[38;2;253;239;231m@\033[38;2;247;229;229m@\033[38;2;232;214;212m&\033[38;2;225;207;204m&\033[38;2;236;218;218m&\033[38;2;229;211;211m&\033[38;2;235;216;221m&\033[38;2;235;216;218m&\033[38;2;242;224;224m&\033[38;2;245;227;227m&\033[38;2;237;219;219m&\033[38;2;233;215;215m&\033[38;2;240;222;222m&\033[38;2;248;230;230m@\033[38;2;233;225;223m&\033[38;2;242;231;232m@\033[38;2;255;253;254m@\033[38;2;178;168;172m*\033[38;2;69;63;65m:\033[38;2;18;16;17m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;6;2;3m \033[38;2;17;8;9m \033[38;2;30;24;24m.\033[38;2;17;13;12m \033[38;2;5;1;2m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;26;6;6m \033[38;2;35;10;13m \033[38;2;25;2;6m \033[38;2;20;0;2m \033[38;2;19;5;5m \033[38;2;17;3;3m \033[38;2;17;3;3m \033[38;2;13;1;1m \033[38;2;12;1;5m \033[38;2;14;1;10m \033[38;2;9;0;7m \033[38;2;11;0;8m \033[38;2;16;3;10m \033[38;2;16;4;8m \033[38;2;16;1;8m \033[38;2;17;1;11m \033[38;2;18;2;12m \033[38;2;17;1;15m \033[38;2;30;13;32m \033[38;2;41;25;44m.\033[38;2;56;45;61m.\033[38;2;73;67;79m:\033[38;2;42;37;52m.\033[38;2;16;15;23m \033[38;2;2;1;6m \033[38;2;1;1;3m \033[38;2;1;1;0m \033[38;2;2;0;1m \033[38;2;5;2;3m \033[38;2;14;3;7m \033[38;2;26;5;5m \033[38;2;141;118;114m=\033[38;2;219;207;193m&\033[38;2;232;212;200m&\033[38;2;240;216;200m&\033[38;2;244;221;205m&\033[38;2;230;218;199m&\033[38;2;253;234;221m@\033[38;2;251;240;231m@\033[38;2;251;248;238m@\033[38;2;254;242;234m@\033[38;2;251;234;228m@\033[38;2;238;213;210m&\033[38;2;214;187;176m#\033[38;2;208;182;169m#\033[38;2;227;197;186m#\033[38;2;238;210;196m&\033[38;2;245;216;200m&\033[38;2;242;210;197m&\033[38;2;231;201;190m&\033[38;2;225;191;181m#\033[38;2;220;185;175m#\033[38;2;221;189;178m#\033[38;2;223;195;179m#\033[38;2;219;191;174m#\033[38;2;201;179;160m#\033[38;2;197;166;156m*\033[38;2;206;171;162m*\033[38;2;188;157;152m*\033[38;2;229;217;207m&\033[38;2;251;251;242m@\033[38;2;246;241;232m@\033[38;2;253;232;228m@\033[38;2;238;217;212m&\033[38;2;224;206;199m&\033[38;2;228;211;203m&\033[38;2;233;213;202m&\033[38;2;227;208;202m&\033[38;2;232;214;212m&\033[38;2;230;211;210m&\033[38;2;231;213;211m&\033[38;2;226;208;208m&\033[38;2;222;204;204m&\033[38;2;229;209;215m&\033[38;2;234;218;219m&\033[38;2;225;214;212m&\033[38;2;228;217;215m&\033[38;2;233;222;220m&\033[38;2;237;222;222m&\033[38;2;238;224;223m&\033[38;2;233;219;218m&\033[38;2;230;221;224m&\033[38;2;230;218;222m&\033[38;2;230;225;230m&\033[38;2;233;228;234m&\033[38;2;43;41;47m.\033[38;2;34;28;38m.\033[38;2;1;0;1m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;5;1;2m \033[38;2;14;8;8m \033[38;2;29;23;23m \033[38;2;8;2;2m \033[38;2;4;0;0m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;47;26;28m.\033[38;2;40;20;21m.\033[38;2;27;5;8m \033[38;2;18;0;1m \033[38;2;12;0;0m \033[38;2;15;1;1m \033[38;2;15;1;1m \033[38;2;12;0;2m \033[38;2;12;0;4m \033[38;2;12;1;7m \033[38;2;11;1;6m \033[38;2;13;2;8m \033[38;2;14;1;8m \033[38;2;14;1;8m \033[38;2;11;0;8m \033[38;2;12;0;8m \033[38;2;16;0;10m \033[38;2;12;0;11m \033[38;2;31;14;31m \033[38;2;53;39;55m.\033[38;2;50;38;52m.\033[38;2;49;41;54m.\033[38;2;39;32;48m.\033[38;2;35;32;41m.\033[38;2;0;0;4m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;4;2;3m \033[38;2;17;8;11m \033[38;2;31;7;9m \033[38;2;171;156;148m*\033[38;2;216;200;187m#\033[38;2;201;181;167m#\033[38;2;225;205;187m&\033[38;2;238;211;194m&\033[38;2;246;220;203m&\033[38;2;225;202;185m#\033[38;2;228;207;191m&\033[38;2;246;220;207m&\033[38;2;243;218;212m&\033[38;2;222;194;186m#\033[38;2;196;165;154m*\033[38;2;200;173;158m*\033[38;2;210;182;168m#\033[38;2;217;186;173m#\033[38;2;236;206;192m&\033[38;2;235;203;191m&\033[38;2;236;204;194m&\033[38;2;232;203;189m&\033[38;2;219;190;176m#\033[38;2;238;209;195m&\033[38;2;251;223;208m&\033[38;2;249;221;210m&\033[38;2;246;218;209m&\033[38;2;249;217;212m&\033[38;2;253;227;217m@\033[38;2;250;230;219m@\033[38;2;248;221;206m&\033[38;2;255;222;210m&\033[38;2;244;216;201m&\033[38;2;240;214;196m&\033[38;2;246;218;206m&\033[38;2;243;214;204m&\033[38;2;235;207;198m&\033[38;2;239;215;207m&\033[38;2;226;209;198m&\033[38;2;227;209;202m&\033[38;2;220;200;199m#\033[38;2;223;203;202m&\033[38;2;220;200;199m#\033[38;2;217;197;196m#\033[38;2;216;196;195m#\033[38;2;222;202;204m&\033[38;2;227;211;209m&\033[38;2;225;211;210m&\033[38;2;223;207;207m&\033[38;2;227;210;212m&\033[38;2;231;215;218m&\033[38;2;231;212;216m&\033[38;2;211;196;199m#\033[38;2;220;215;209m&\033[38;2;221;215;212m&\033[38;2;224;216;220m&\033[38;2;214;209;213m&\033[38;2;70;65;72m:\033[38;2;38;35;43m.\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;4;0;1m \033[38;2;10;1;2m \033[38;2;7;1;1m \033[38;2;14;8;8m \033[38;2;1;1;1m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;44;30;30m.\033[38;2;38;24;24m.\033[38;2;24;8;9m \033[38;2;17;1;2m \033[38;2;17;5;7m \033[38;2;26;14;16m \033[38;2;39;27;29m.\033[38;2;22;7;10m \033[38;2;16;1;4m \033[38;2;9;0;0m \033[38;2;9;0;1m \033[38;2;11;0;4m \033[38;2;13;0;9m \033[38;2;14;1;10m \033[38;2;15;4;12m \033[38;2;13;0;9m \033[38;2;14;1;10m \033[38;2;23;7;9m \033[38;2;91;76;86m-\033[38;2;87;76;84m-\033[38;2;87;75;85m-\033[38;2;63;52;68m:\033[38;2;49;40;57m.\033[38;2;26;20;32m \033[38;2;1;0;11m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;2;0;3m \033[38;2;17;9;10m \033[38;2;30;7;9m \033[38;2;192;181;173m#\033[38;2;219;204;195m#\033[38;2;182;165;149m*\033[38;2;196;175;159m*\033[38;2;211;185;168m#\033[38;2;223;197;184m#\033[38;2;229;203;190m&\033[38;2;234;208;193m&\033[38;2;224;196;182m#\033[38;2;206;173;154m*\033[38;2;174;132;111m+\033[38;2;167;131;107m+\033[38;2;207;171;154m*\033[38;2;208;173;154m*\033[38;2;176;143;124m+\033[38;2;167;129;112m+\033[38;2;169;141;116m+\033[38;2;234;194;178m#\033[38;2;235;204;184m&\033[38;2;253;223;206m&\033[38;2;247;220;204m&\033[38;2;239;211;199m&\033[38;2;248;222;207m&\033[38;2;254;233;216m@\033[38;2;234;202;191m&\033[38;2;240;210;198m&\033[38;2;242;212;201m&\033[38;2;241;214;203m&\033[38;2;248;221;210m&\033[38;2;251;224;214m&\033[38;2;247;224;210m&\033[38;2;244;223;206m&\033[38;2;240;218;204m&\033[38;2;230;211;197m&\033[38;2;209;190;176m#\033[38;2;200;182;171m#\033[38;2;196;179;169m#\033[38;2;193;174;168m*\033[38;2;201;182;176m#\033[38;2;206;187;181m#\033[38;2;203;184;178m#\033[38;2;204;185;179m#\033[38;2;203;184;180m#\033[38;2;210;191;187m#\033[38;2;208;189;185m#\033[38;2;207;189;189m#\033[38;2;205;187;187m#\033[38;2;218;199;203m#\033[38;2;227;206;211m&\033[38;2;216;199;204m#\033[38;2;206;201;205m#\033[38;2;210;205;202m#\033[38;2;213;206;215m&\033[38;2;232;221;227m&\033[38;2;104;98;111m-\033[38;2;33;30;40m.\033[38;2;5;5;3m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;0;1m \033[38;2;10;1;2m \033[38;2;9;0;1m \033[38;2;9;0;1m \033[38;2;3;1;2m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;26;12;12m \033[38;2;28;14;14m \033[38;2;14;0;0m \033[38;2;26;6;8m \033[38;2;13;1;3m \033[38;2;12;0;2m \033[38;2;14;1;3m \033[38;2;17;2;5m \033[38;2;16;1;4m \033[38;2;14;0;3m \033[38;2;8;0;1m \033[38;2;10;1;5m \033[38;2;13;1;3m \033[38;2;12;0;2m \033[38;2;13;1;6m \033[38;2;16;1;6m \033[38;2;20;3;9m \033[38;2;20;1;3m \033[38;2;22;5;15m \033[38;2;62;46;57m:\033[38;2;64;48;59m:\033[38;2;38;24;41m.\033[38;2;39;24;45m.\033[38;2;24;11;31m \033[38;2;8;2;15m \033[38;2;1;1;6m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;2;0;3m \033[38;2;16;7;8m \033[38;2;26;3;7m \033[38;2;187;175;170m*\033[38;2;210;198;186m#\033[38;2;170;146;139m+\033[38;2;153;121;110m=\033[38;2;154;121;106m=\033[38;2;177;147;134m+\033[38;2;216;186;179m#\033[38;2;212;185;176m#\033[38;2;226;205;192m&\033[38;2;251;222;204m&\033[38;2;189;151;132m*\033[38;2;113;61;38m:\033[38;2;132;81;51m-\033[38;2;145;82;64m-\033[38;2;93;17;9m.\033[38;2;104;2;2m.\033[38;2;104;27;14m.\033[38;2;157;125;100m+\033[38;2;197;159;144m*\033[38;2;245;214;199m&\033[38;2;248;223;209m&\033[38;2;236;214;201m&\033[38;2;237;210;196m&\033[38;2;242;213;200m&\033[38;2;230;200;189m&\033[38;2;238;210;198m&\033[38;2;239;212;199m&\033[38;2;234;207;196m&\033[38;2;234;207;196m&\033[38;2;228;204;194m&\033[38;2;216;194;180m#\033[38;2;209;190;173m#\033[38;2;206;184;170m#\033[38;2;194;175;161m*\033[38;2;190;171;158m*\033[38;2;179;160;149m*\033[38;2;174;157;147m*\033[38;2;181;162;156m*\033[38;2;198;179;173m#\033[38;2;202;183;177m#\033[38;2;208;189;183m#\033[38;2;214;195;189m#\033[38;2;205;186;179m#\033[38;2;195;176;169m*\033[38;2;196;177;170m#\033[38;2;190;171;164m*\033[38;2;188;168;167m*\033[38;2;195;175;176m*\033[38;2;205;183;186m#\033[38;2;203;184;188m#\033[38;2;200;189;197m#\033[38;2;215;206;209m&\033[38;2;216;207;218m&\033[38;2;217;212;216m&\033[38;2;143;137;150m+\033[38;2;28;17;33m \033[38;2;10;8;11m \033[38;2;0;1;5m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;5;1;2m \033[38;2;9;5;6m \033[38;2;7;3;4m \033[38;2;5;1;2m \033[38;2;2;0;1m \033[38;2;1;1;3m \033[0m");
        $display("\033[38;2;26;6;8m \033[38;2;12;0;0m \033[38;2;9;3;0m \033[38;2;17;1;2m \033[38;2;10;0;1m \033[38;2;10;0;1m \033[38;2;16;1;4m \033[38;2;34;19;22m \033[38;2;17;5;7m \033[38;2;10;0;1m \033[38;2;9;0;1m \033[38;2;16;4;8m \033[38;2;28;13;16m \033[38;2;17;5;7m \033[38;2;14;2;6m \033[38;2;21;4;10m \033[38;2;22;3;9m \033[38;2;40;19;28m.\033[38;2;21;4;14m \033[38;2;23;7;19m \033[38;2;53;41;51m.\033[38;2;44;33;49m.\033[38;2;28;17;33m \033[38;2;24;12;32m \033[38;2;6;0;12m \033[38;2;1;0;5m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;5;2;1m \033[38;2;15;6;6m \033[38;2;31;6;6m \033[38;2;184;174;169m*\033[38;2;215;204;200m#\033[38;2;164;145;139m+\033[38;2;149;120;116m=\033[38;2;146;115;111m=\033[38;2;174;144;142m+\033[38;2;193;160;155m*\033[38;2;213;182;177m#\033[38;2;229;202;193m&\033[38;2;226;199;190m#\033[38;2;249;221;209m&\033[38;2;209;172;158m*\033[38;2;122;57;44m:\033[38;2;122;51;33m:\033[38;2;177;130;114m+\033[38;2;233;200;188m&\033[38;2;249;217;205m&\033[38;2;253;232;227m@\033[38;2;253;230;216m@\033[38;2;242;217;204m&\033[38;2;252;229;213m@\033[38;2;241;213;199m&\033[38;2;233;207;189m&\033[38;2;225;199;184m#\033[38;2;217;189;175m#\033[38;2;222;196;181m#\033[38;2;214;191;175m#\033[38;2;210;187;171m#\033[38;2;205;182;168m#\033[38;2;186;164;150m*\033[38;2;171;150;133m+\033[38;2;160;141;124m+\033[38;2;135;117;95m=\033[38;2;132;114;94m=\033[38;2;137;118;103m=\033[38;2;151;132;115m+\033[38;2;166;148;135m+\033[38;2;192;174;164m*\033[38;2;193;175;165m*\033[38;2;195;177;167m*\033[38;2;202;184;174m#\033[38;2;189;171;161m*\033[38;2;200;181;174m#\033[38;2;206;187;180m#\033[38;2;204;185;178m#\033[38;2;205;188;180m#\033[38;2;205;188;181m#\033[38;2;208;191;185m#\033[38;2;207;186;185m#\033[38;2;193;172;177m*\033[38;2;186;175;181m*\033[38;2;189;178;186m#\033[38;2;208;197;211m#\033[38;2;195;187;200m#\033[38;2;86;78;99m-\033[38;2;20;10;31m \033[38;2;7;6;10m \033[38;2;3;1;4m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;5;1;0m \033[38;2;6;2;3m \033[38;2;5;1;1m \033[38;2;5;1;2m \033[38;2;1;0;0m \033[38;2;1;1;3m \033[0m");
        $display("\033[38;2;16;0;1m \033[38;2;20;0;2m \033[38;2;31;8;11m \033[38;2;43;20;24m.\033[38;2;24;5;9m \033[38;2;28;9;13m \033[38;2;26;7;11m \033[38;2;23;6;7m \033[38;2;24;8;9m \033[38;2;20;4;7m \033[38;2;12;1;2m \033[38;2;11;1;2m \033[38;2;12;0;2m \033[38;2;20;7;10m \033[38;2;15;3;5m \033[38;2;12;2;3m \033[38;2;17;2;5m \033[38;2;29;14;21m \033[38;2;42;27;37m.\033[38;2;59;49;57m:\033[38;2;56;49;57m:\033[38;2;44;38;52m.\033[38;2;28;21;37m \033[38;2;35;27;48m.\033[38;2;7;0;16m \033[38;2;9;4;15m \033[38;2;3;0;6m \033[38;2;5;1;2m \033[38;2;10;4;4m \033[38;2;15;0;3m \033[38;2;33;2;2m \033[38;2;157;148;141m+\033[38;2;184;169;166m*\033[38;2;143;124;117m=\033[38;2;143;124;117m=\033[38;2;151;124;118m+\033[38;2;135;116;101m=\033[38;2;146;122;112m=\033[38;2;157;131;118m+\033[38;2;179;151;142m*\033[38;2;196;169;162m*\033[38;2;185;157;151m*\033[38;2;173;143;138m+\033[38;2;164;123;122m+\033[38;2;131;85;83m-\033[38;2;166;125;121m+\033[38;2;179;133;130m+\033[38;2;183;144;139m+\033[38;2;199;166;157m*\033[38;2;200;174;162m*\033[38;2;208;186;172m#\033[38;2;205;178;165m#\033[38;2;199;168;157m*\033[38;2;201;172;164m*\033[38;2;202;177;170m#\033[38;2;214;185;174m#\033[38;2;203;177;164m#\033[38;2;200;181;167m#\033[38;2;205;186;172m#\033[38;2;188;169;155m*\033[38;2;157;135;121m+\033[38;2;138;119;105m=\033[38;2;157;138;124m+\033[38;2;175;153;142m*\033[38;2;184;162;151m*\033[38;2;198;176;165m*\033[38;2;187;165;154m*\033[38;2;197;175;164m*\033[38;2;209;192;184m#\033[38;2;207;188;182m#\033[38;2;199;180;173m#\033[38;2;199;180;173m#\033[38;2;207;188;180m#\033[38;2;210;192;182m#\033[38;2;211;193;183m#\033[38;2;207;189;179m#\033[38;2;213;196;188m#\033[38;2;215;200;193m#\033[38;2;213;198;197m#\033[38;2;223;205;208m&\033[38;2;225;208;214m&\033[38;2;220;211;210m&\033[38;2;221;213;219m&\033[38;2;211;203;213m#\033[38;2;203;197;207m#\033[38;2;121;115;127m=\033[38;2;31;23;36m.\033[38;2;19;18;23m \033[38;2;2;0;5m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;3;1;2m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[0m");
        $display("\033[38;2;18;0;2m \033[38;2;19;0;2m \033[38;2;24;2;5m \033[38;2;30;8;9m \033[38;2;25;9;10m \033[38;2;18;2;3m \033[38;2;15;0;0m \033[38;2;13;1;3m \033[38;2;13;1;3m \033[38;2;11;1;2m \033[38;2;5;0;0m \033[38;2;14;4;5m \033[38;2;16;6;7m \033[38;2;10;0;1m \033[38;2;12;0;2m \033[38;2;10;0;0m \033[38;2;29;14;17m \033[38;2;40;27;37m.\033[38;2;68;56;64m:\033[38;2;63;55;62m:\033[38;2;51;46;52m.\033[38;2;45;34;48m.\033[38;2;27;19;39m \033[38;2;26;17;34m \033[38;2;15;6;23m \033[38;2;39;28;42m.\033[38;2;32;19;29m \033[38;2;10;1;4m \033[38;2;12;0;2m \033[38;2;16;1;4m \033[38;2;43;9;10m \033[38;2;123;107;102m=\033[38;2;209;191;191m#\033[38;2;175;157;147m*\033[38;2;142;122;115m=\033[38;2;159;137;128m+\033[38;2;134;109;94m=\033[38;2;137;114;96m=\033[38;2;138;112;99m=\033[38;2;162;134;126m+\033[38;2;153;124;116m+\033[38;2;103;63;63m:\033[38;2;92;48;48m:\033[38;2;70;18;19m.\033[38;2;68;1;3m \033[38;2;105;40;41m:\033[38;2;109;59;55m:\033[38;2;157;119;110m=\033[38;2;176;146;136m+\033[38;2;193;166;159m*\033[38;2;188;157;152m*\033[38;2;189;159;153m*\033[38;2;184;162;154m*\033[38;2;185;162;151m*\033[38;2;189;162;150m*\033[38;2;183;153;145m*\033[38;2;179;151;143m*\033[38;2;182;155;146m*\033[38;2;185;163;152m*\033[38;2;172;150;137m+\033[38;2;156;135;121m+\033[38;2;152;130;117m+\033[38;2;167;145;132m+\033[38;2;191;173;163m*\033[38;2;195;176;167m*\033[38;2;184;166;156m*\033[38;2;179;159;148m*\033[38;2;181;161;151m*\033[38;2;202;185;175m#\033[38;2;217;198;188m#\033[38;2;196;178;168m#\033[38;2;210;192;182m#\033[38;2;205;187;177m#\033[38;2;206;188;178m#\033[38;2;203;185;175m#\033[38;2;205;187;177m#\033[38;2;213;196;188m#\033[38;2;221;203;198m&\033[38;2;223;207;207m&\033[38;2;229;213;216m&\033[38;2;226;210;213m&\033[38;2;217;207;207m&\033[38;2;221;212;215m&\033[38;2;206;198;206m#\033[38;2;197;191;203m#\033[38;2;191;185;197m#\033[38;2;85;75;89m-\033[38;2;9;8;14m \033[38;2;2;1;6m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;2;1;2m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;28;8;10m \033[38;2;22;1;3m \033[38;2;26;4;6m \033[38;2;43;21;22m.\033[38;2;26;7;9m \033[38;2;15;0;0m \033[38;2;13;0;0m \033[38;2;13;0;2m \033[38;2;15;2;4m \033[38;2;13;1;3m \033[38;2;9;0;1m \033[38;2;11;0;2m \033[38;2;17;2;5m \033[38;2;14;0;2m \033[38;2;21;6;9m \033[38;2;14;0;2m \033[38;2;13;1;3m \033[38;2;16;0;9m \033[38;2;38;22;32m.\033[38;2;58;41;51m.\033[38;2;56;45;53m.\033[38;2;49;41;54m.\033[38;2;50;39;57m.\033[38;2;10;2;14m \033[38;2;10;3;10m \033[38;2;14;4;12m \033[38;2;45;33;41m.\033[38;2;15;3;7m \033[38;2;20;5;8m \033[38;2;19;2;5m \033[38;2;29;1;0m \033[38;2;125;115;109m=\033[38;2;188;172;173m*\033[38;2;183;166;159m*\033[38;2;184;166;162m*\033[38;2;178;157;149m*\033[38;2;164;147;129m+\033[38;2;142;123;105m=\033[38;2;99;71;60m-\033[38;2;79;29;30m.\033[38;2;67;18;21m.\033[38;2;35;1;0m \033[38;2;30;0;0m \033[38;2;31;1;1m \033[38;2;38;1;0m \033[38;2;42;2;5m \033[38;2;39;0;1m \033[38;2;37;0;1m \033[38;2;43;1;1m \033[38;2;58;1;3m \033[38;2;84;29;29m.\033[38;2;99;52;49m:\033[38;2;146;116;107m=\033[38;2;157;131;124m+\033[38;2;159;133;128m+\033[38;2;170;144;137m+\033[38;2;172;145;138m+\033[38;2;162;133;127m+\033[38;2;148;120;112m=\033[38;2;132;104;93m=\033[38;2;112;85;71m-\033[38;2;96;70;53m:\033[38;2;120;93;77m-\033[38;2;140;120;102m=\033[38;2;141;120;107m=\033[38;2;171;149;141m+\033[38;2;190;170;159m*\033[38;2;200;180;169m#\033[38;2;189;171;157m*\033[38;2;179;160;146m*\033[38;2;194;176;162m*\033[38;2;200;182;168m#\033[38;2;191;173;159m*\033[38;2;202;184;170m#\033[38;2;217;199;185m#\033[38;2;220;202;188m#\033[38;2;223;206;198m&\033[38;2;220;203;197m#\033[38;2;217;202;202m#\033[38;2;226;210;213m&\033[38;2;223;207;210m&\033[38;2;217;208;211m&\033[38;2;220;208;216m&\033[38;2;223;213;224m&\033[38;2;206;200;212m#\033[38;2;182;178;190m*\033[38;2;91;85;93m-\033[38;2;30;27;33m.\033[38;2;4;1;4m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;1;2m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;3;0;2m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;37;16;17m \033[38;2;37;17;17m \033[38;2;51;29;31m.\033[38;2;60;38;40m.\033[38;2;34;20;20m \033[38;2;15;1;1m \033[38;2;15;1;1m \033[38;2;15;0;3m \033[38;2;18;3;6m \033[38;2;17;4;6m \033[38;2;12;1;2m \033[38;2;12;0;2m \033[38;2;13;0;2m \033[38;2;17;1;4m \033[38;2;16;1;3m \033[38;2;24;7;10m \033[38;2;30;11;15m \033[38;2;43;26;32m.\033[38;2;53;40;47m.\033[38;2;69;56;65m:\033[38;2;48;38;46m.\033[38;2;45;36;47m.\033[38;2;28;22;36m \033[38;2;9;1;17m \033[38;2;17;9;23m \033[38;2;46;34;48m.\033[38;2;25;13;23m \033[38;2;21;7;17m \033[38;2;11;1;5m \033[38;2;29;15;19m \033[38;2;26;5;5m \033[38;2;155;146;141m+\033[38;2;202;195;184m#\033[38;2;184;172;158m*\033[38;2;191;168;155m*\033[38;2;191;172;155m*\033[38;2;175;169;143m*\033[38;2;178;166;143m*\033[38;2;151;131;113m+\033[38;2;126;101;87m=\033[38;2;85;46;44m:\033[38;2;78;29;32m.\033[38;2;53;4;5m \033[38;2;82;40;41m:\033[38;2;115;78;79m-\033[38;2;118;86;90m-\033[38;2;135;97;103m=\033[38;2;129;89;95m-\033[38;2;97;53;58m:\033[38;2;76;35;30m.\033[38;2;44;0;0m \033[38;2;49;0;1m \033[38;2;55;0;1m \033[38;2;55;2;1m \033[38;2;73;14;13m.\033[38;2;104;50;41m:\033[38;2;78;20;12m.\033[38;2;66;10;3m.\033[38;2;69;15;3m.\033[38;2;94;53;42m:\033[38;2;101;68;61m:\033[38;2;122;97;91m=\033[38;2;135;112;100m=\033[38;2;152;126;113m+\033[38;2;149;125;111m+\033[38;2;162;139;123m+\033[38;2;162;134;117m+\033[38;2;160;128;112m+\033[38;2;174;147;133m+\033[38;2;192;165;153m*\033[38;2;192;165;154m*\033[38;2;183;159;151m*\033[38;2;202;179;171m#\033[38;2;212;192;188m#\033[38;2;207;190;182m#\033[38;2;202;189;177m#\033[38;2;208;194;187m#\033[38;2;206;194;190m#\033[38;2;203;192;188m#\033[38;2;200;189;191m#\033[38;2;207;196;197m#\033[38;2;190;180;188m#\033[38;2;199;191;205m#\033[38;2;200;192;207m#\033[38;2;183;180;190m#\033[38;2;164;163;168m*\033[38;2;55;53;64m:\033[38;2;23;22;29m \033[38;2;4;3;9m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[0m");
        $display("\033[38;2;24;4;9m \033[38;2;31;11;12m \033[38;2;28;8;9m \033[38;2;22;0;2m \033[38;2;19;0;3m \033[38;2;22;3;6m \033[38;2;19;5;6m \033[38;2;16;1;4m \033[38;2;15;0;3m \033[38;2;12;0;2m \033[38;2;8;0;0m \033[38;2;11;0;2m \033[38;2;12;0;2m \033[38;2;17;1;2m \033[38;2;16;1;4m \033[38;2;35;19;22m \033[38;2;50;35;38m.\033[38;2;40;25;30m.\033[38;2;44;28;36m.\033[38;2;51;37;45m.\033[38;2;48;40;48m.\033[38;2;44;39;46m.\033[38;2;41;33;46m.\033[38;2;20;11;28m \033[38;2;10;2;17m \033[38;2;33;25;36m.\033[38;2;35;24;33m.\033[38;2;8;1;6m \033[38;2;5;3;1m \033[38;2;10;1;2m \033[38;2;36;14;16m \033[38;2;156;136;135m+\033[38;2;181;171;162m*\033[38;2;184;170;161m*\033[38;2;193;172;162m*\033[38;2;186;169;155m*\033[38;2;181;168;150m*\033[38;2;196;178;166m#\033[38;2;171;153;141m*\033[38;2;139;115;105m=\033[38;2;127;99;94m=\033[38;2;158;127;123m+\033[38;2;153;126;117m+\033[38;2;171;142;134m+\033[38;2;172;147;139m+\033[38;2;160;132;122m+\033[38;2;156;123;115m+\033[38;2;164;131;121m+\033[38;2;182;153;144m*\033[38;2;166;137;129m+\033[38;2;157;129;124m+\033[38;2;144;116;111m=\033[38;2;156;125;127m+\033[38;2;151;124;123m+\033[38;2;153;126;128m+\033[38;2;136;109;102m=\033[38;2;124;98;92m=\033[38;2;126;96;92m=\033[38;2;128;102;91m=\033[38;2;147;127;118m+\033[38;2;150;130;123m+\033[38;2;172;154;144m*\033[38;2;185;167;155m*\033[38;2;200;182;170m#\033[38;2;202;182;171m#\033[38;2;210;188;177m#\033[38;2;222;195;183m#\033[38;2;216;187;173m#\033[38;2;211;185;170m#\033[38;2;195;169;155m*\033[38;2;197;171;161m*\033[38;2;198;176;165m*\033[38;2;201;181;170m#\033[38;2;201;176;169m#\033[38;2;203;187;177m#\033[38;2;203;191;179m#\033[38;2;197;183;175m#\033[38;2;195;184;180m#\033[38;2;197;187;184m#\033[38;2;194;183;187m#\033[38;2;199;188;194m#\033[38;2;191;184;191m#\033[38;2;196;188;199m#\033[38;2;186;180;193m#\033[38;2;201;198;208m#\033[38;2;170;169;177m*\033[38;2;27;26;34m.\033[38;2;20;19;25m \033[38;2;2;1;6m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[0m");
        $display("\033[38;2;20;1;3m \033[38;2;24;4;3m \033[38;2;39;18;20m \033[38;2;34;12;14m \033[38;2;20;2;6m \033[38;2;23;4;8m \033[38;2;12;1;2m \033[38;2;11;1;0m \033[38;2;12;0;2m \033[38;2;16;1;4m \033[38;2;9;0;2m \033[38;2;13;0;4m \033[38;2;14;1;0m \033[38;2;16;0;1m \033[38;2;23;4;6m \033[38;2;17;1;2m \033[38;2;45;29;32m.\033[38;2;41;27;28m.\033[38;2;43;28;36m.\033[38;2;52;38;48m.\033[38;2;42;35;42m.\033[38;2;39;32;40m.\033[38;2;32;26;40m.\033[38;2;12;4;20m \033[38;2;37;24;42m.\033[38;2;33;25;33m.\033[38;2;19;7;15m \033[38;2;13;0;9m \033[38;2;10;0;1m \033[38;2;10;0;1m \033[38;2;22;2;4m \033[38;2;52;27;30m.\033[38;2;157;143;140m+\033[38;2;175;161;157m*\033[38;2;185;167;158m*\033[38;2;182;165;155m*\033[38;2;168;152;139m+\033[38;2;179;159;148m*\033[38;2;163;144;130m+\033[38;2;149;125;113m+\033[38;2;117;94;76m-\033[38;2;122;93;77m-\033[38;2;145;118;102m=\033[38;2;177;154;140m*\033[38;2;160;136;124m+\033[38;2;156;128;117m+\033[38;2;140;106;96m=\033[38;2;134;102;90m=\033[38;2;147;115;104m=\033[38;2;145;115;106m=\033[38;2;151;123;119m+\033[38;2;154;130;122m+\033[38;2;179;158;153m*\033[38;2;174;153;151m*\033[38;2;143;121;123m=\033[38;2;126;105;104m=\033[38;2;130;108;109m=\033[38;2;127;106;103m=\033[38;2;120;100;86m=\033[38;2;138;111;97m=\033[38;2;133;109;92m=\033[38;2;158;138;123m+\033[38;2;165;148;135m+\033[38;2;183;162;149m*\033[38;2;180;158;145m*\033[38;2;181;158;144m*\033[38;2;191;164;150m*\033[38;2;198;170;156m*\033[38;2;222;196;182m#\033[38;2;214;188;171m#\033[38;2;210;184;166m#\033[38;2;181;157;145m*\033[38;2;190;171;157m*\033[38;2;186;166;157m*\033[38;2;175;158;150m*\033[38;2;172;159;146m*\033[38;2;177;164;156m*\033[38;2;178;167;165m*\033[38;2;189;182;175m#\033[38;2;185;176;176m*\033[38;2;186;175;181m*\033[38;2;194;188;195m#\033[38;2;191;181;191m#\033[38;2;172;166;178m*\033[38;2;152;150;165m+\033[38;2;65;63;74m:\033[38;2;25;24;30m \033[38;2;6;6;8m \033[38;2;0;0;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;18;2;5m \033[38;2;20;1;3m \033[38;2;35;17;17m \033[38;2;34;14;15m \033[38;2;22;6;9m \033[38;2;11;0;1m \033[38;2;11;0;1m \033[38;2;11;1;0m \033[38;2;11;0;1m \033[38;2;15;0;3m \033[38;2;13;3;4m \033[38;2;13;0;4m \033[38;2;21;5;6m \033[38;2;25;6;7m \033[38;2;21;2;4m \033[38;2;16;0;1m \033[38;2;51;35;38m.\033[38;2;43;28;31m.\033[38;2;45;30;37m.\033[38;2;53;39;48m.\033[38;2;28;20;28m \033[38;2;38;31;39m.\033[38;2;45;37;52m.\033[38;2;21;12;29m \033[38;2;29;21;36m \033[38;2;16;5;21m \033[38;2;12;0;11m \033[38;2;15;2;10m \033[38;2;13;3;4m \033[38;2;8;0;0m \033[38;2;12;2;3m \033[38;2;25;6;8m \033[38;2;124;108;108m=\033[38;2;180;166;164m*\033[38;2;154;135;129m+\033[38;2;133;113;107m=\033[38;2;178;158;151m*\033[38;2;179;159;152m*\033[38;2;161;141;131m+\033[38;2;142;118;108m=\033[38;2;127;104;90m=\033[38;2;110;91;76m-\033[38;2;105;83;70m-\033[38;2;125;105;95m=\033[38;2;121;101;94m=\033[38;2;149;122;115m=\033[38;2;142;112;105m=\033[38;2;145;115;106m=\033[38;2;138;109;101m=\033[38;2;124;98;83m=\033[38;2;125;98;91m=\033[38;2;133;110;100m=\033[38;2;121;100;94m=\033[38;2;122;103;99m=\033[38;2;90;72;66m:\033[38;2;78;60;55m:\033[38;2;81;61;60m:\033[38;2;88;69;63m:\033[38;2;86;67;53m:\033[38;2;126;105;88m=\033[38;2;165;150;129m+\033[38;2;202;186;170m#\033[38;2;198;183;170m#\033[38;2;215;197;185m#\033[38;2;195;175;164m*\033[38;2;195;173;161m*\033[38;2;197;171;158m*\033[38;2;197;170;158m*\033[38;2;184;158;143m*\033[38;2;185;159;144m*\033[38;2;189;164;147m*\033[38;2;178;157;143m*\033[38;2;178;160;146m*\033[38;2;177;158;141m*\033[38;2;173;156;144m*\033[38;2;182;170;157m*\033[38;2;185;172;164m*\033[38;2;182;171;169m*\033[38;2;168;161;158m*\033[38;2;171;165;169m*\033[38;2;170;160;167m*\033[38;2;167;160;167m*\033[38;2;154;144;153m+\033[38;2;99;92;107m-\033[38;2;94;91;112m-\033[38;2;51;47;63m.\033[38;2;4;1;17m \033[38;2;10;9;15m \033[38;2;3;2;7m \033[38;2;0;0;4m \033[38;2;1;1;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;29;14;19m \033[38;2;20;5;10m \033[38;2;16;1;4m \033[38;2;16;2;4m \033[38;2;18;4;4m \033[38;2;15;3;5m \033[38;2;12;0;4m \033[38;2;12;2;3m \033[38;2;9;0;0m \033[38;2;16;4;4m \033[38;2;9;2;1m \033[38;2;9;1;0m \033[38;2;13;1;3m \033[38;2;13;1;3m \033[38;2;15;0;3m \033[38;2;41;26;29m.\033[38;2;58;41;46m.\033[38;2;33;14;18m \033[38;2;21;5;11m \033[38;2;53;40;46m.\033[38;2;52;42;50m.\033[38;2;48;41;49m.\033[38;2;37;30;38m.\033[38;2;18;10;23m \033[38;2;12;4;19m \033[38;2;31;19;33m \033[38;2;27;15;25m \033[38;2;15;4;10m \033[38;2;12;6;10m \033[38;2;3;1;4m \033[38;2;5;1;2m \033[38;2;18;6;6m \033[38;2;19;5;5m \033[38;2;143;129;128m+\033[38;2;174;160;159m*\033[38;2;166;152;151m*\033[38;2;165;150;145m+\033[38;2;156;137;130m+\033[38;2;144;127;117m+\033[38;2;156;139;129m+\033[38;2;147;130;123m+\033[38;2;138;119;113m=\033[38;2;114;97;90m-\033[38;2;108;92;82m-\033[38;2;96;78;68m-\033[38;2;83;58;53m:\033[38;2;69;44;39m.\033[38;2;69;42;38m.\033[38;2;86;59;53m:\033[38;2;67;42;35m.\033[38;2;66;42;36m.\033[38;2;66;38;34m.\033[38;2;39;11;12m \033[38;2;34;13;8m \033[38;2;28;7;6m \033[38;2;26;1;0m \033[38;2;30;6;4m \033[38;2;50;29;26m.\033[38;2;85;64;63m:\033[38;2;131;111;110m=\033[38;2;130;109;106m=\033[38;2;125;104;99m=\033[38;2;128;99;97m=\033[38;2;132;102;100m=\033[38;2;135;105;103m=\033[38;2;140;110;108m=\033[38;2;138;100;101m=\033[38;2;135;92;94m=\033[38;2;115;85;77m-\033[38;2;125;97;88m=\033[38;2;138;110;101m=\033[38;2;143;123;109m=\033[38;2;148;133;118m+\033[38;2;138;126;112m=\033[38;2;129;114;97m=\033[38;2;115;98;78m-\033[38;2;117;105;85m=\033[38;2;146;135;121m+\033[38;2;132;121;117m=\033[38;2;149;137;139m+\033[38;2;141;128;137m+\033[38;2;123;121;132m=\033[38;2;112;110;121m=\033[38;2;146;144;155m+\033[38;2;151;150;158m+\033[38;2;155;154;160m+\033[38;2;109;107;113m=\033[38;2;60;59;64m:\033[38;2;8;7;12m \033[38;2;1;0;2m \033[38;2;2;0;1m \033[38;2;1;0;0m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;26;16;22m \033[38;2;17;8;13m \033[38;2;9;0;3m \033[38;2;11;2;5m \033[38;2;7;3;4m \033[38;2;4;0;1m \033[38;2;5;1;2m \033[38;2;4;0;1m \033[38;2;6;2;3m \033[38;2;6;2;3m \033[38;2;3;1;2m \033[38;2;0;0;0m \033[38;2;3;0;0m \033[38;2;4;0;0m \033[38;2;4;0;1m \033[38;2;4;0;1m \033[38;2;9;3;5m \033[38;2;5;0;1m \033[38;2;5;2;3m \033[38;2;5;1;4m \033[38;2;4;1;5m \033[38;2;4;2;7m \033[38;2;1;0;6m \033[38;2;1;1;3m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;4;3;4m \033[38;2;5;5;7m \033[38;2;13;7;11m \033[38;2;16;1;3m \033[38;2;19;9;10m \033[38;2;24;15;16m \033[38;2;54;42;44m.\033[38;2;51;41;42m.\033[38;2;66;61;61m:\033[38;2;66;63;62m:\033[38;2;65;62;61m:\033[38;2;65;62;61m:\033[38;2;66;61;63m:\033[38;2;66;60;64m:\033[38;2;64;60;64m:\033[38;2;62;61;64m:\033[38;2;57;55;58m:\033[38;2;56;47;50m.\033[38;2;62;47;52m:\033[38;2;54;42;45m.\033[38;2;48;36;38m.\033[38;2;44;31;33m.\033[38;2;42;33;35m.\033[38;2;39;32;34m.\033[38;2;34;34;36m.\033[38;2;37;35;36m.\033[38;2;36;33;34m.\033[38;2;34;29;33m.\033[38;2;35;30;34m.\033[38;2;17;15;18m \033[38;2;40;29;33m.\033[38;2;43;33;34m.\033[38;2;43;33;31m.\033[38;2;45;33;33m.\033[38;2;44;35;37m.\033[38;2;41;30;31m.\033[38;2;42;28;28m.\033[38;2;40;24;25m.\033[38;2;35;16;15m \033[38;2;30;5;7m \033[38;2;42;20;22m.\033[38;2;37;11;10m \033[38;2;34;5;3m \033[38;2;32;2;1m \033[38;2;35;1;1m \033[38;2;33;0;0m \033[38;2;32;0;0m \033[38;2;32;2;2m \033[38;2;41;11;9m \033[38;2;43;17;16m \033[38;2;30;4;2m \033[38;2;30;6;6m \033[38;2;22;0;3m \033[38;2;18;1;20m \033[38;2;27;10;29m \033[38;2;15;3;18m \033[38;2;6;1;7m \033[38;2;23;21;26m \033[38;2;18;16;17m \033[38;2;6;4;5m \033[38;2;4;2;3m \033[38;2;2;0;1m \033[38;2;1;1;1m \033[38;2;1;0;0m \033[38;2;4;2;3m \033[38;2;4;2;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;0;1m \033[38;2;2;0;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;1;1;3m \033[38;2;1;1;2m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;1;0m \033[38;2;0;1;0m \033[38;2;0;0;0m \033[38;2;2;0;3m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[38;2;1;0;6m \033[38;2;4;3;8m \033[38;2;12;11;13m \033[38;2;34;28;35m.\033[38;2;58;51;61m:\033[38;2;79;72;79m:\033[38;2;72;62;72m:\033[38;2;52;40;54m.\033[38;2;137;127;130m+\033[38;2;219;209;212m&\033[38;2;229;225;226m&\033[38;2;240;239;239m@\033[38;2;246;243;243m@\033[38;2;248;247;247m@\033[38;2;250;248;249m@\033[38;2;247;247;247m@\033[38;2;250;249;249m@\033[38;2;252;248;247m@\033[38;2;251;248;249m@\033[38;2;253;250;253m@\033[38;2;254;252;254m@\033[38;2;254;253;254m@\033[38;2;253;253;253m@\033[38;2;254;251;252m@\033[38;2;252;249;250m@\033[38;2;252;249;250m@\033[38;2;252;249;252m@\033[38;2;248;249;246m@\033[38;2;249;246;247m@\033[38;2;247;245;246m@\033[38;2;247;245;246m@\033[38;2;248;245;246m@\033[38;2;248;245;246m@\033[38;2;248;243;237m@\033[38;2;247;241;238m@\033[38;2;249;242;244m@\033[38;2;242;234;232m@\033[38;2;238;224;222m&\033[38;2;231;218;214m&\033[38;2;227;216;208m&\033[38;2;230;220;209m&\033[38;2;230;219;207m&\033[38;2;229;215;204m&\033[38;2;222;207;197m&\033[38;2;222;204;196m&\033[38;2;222;199;193m#\033[38;2;215;185;189m#\033[38;2;220;191;195m#\033[38;2;230;204;207m&\033[38;2;225;203;201m&\033[38;2;221;198;199m#\033[38;2;209;194;192m#\033[38;2;203;187;184m#\033[38;2;195;179;175m#\033[38;2;194;181;178m#\033[38;2;184;174;173m*\033[38;2;180;174;173m*\033[38;2;183;179;178m*\033[38;2;177;172;172m*\033[38;2;144;134;142m+\033[38;2;106;96;104m-\033[38;2;96;85;93m-\033[38;2;62;49;57m:\033[38;2;36;23;29m.\033[38;2;63;53;56m:\033[38;2;77;71;73m:\033[38;2;89;81;84m-\033[38;2;98;84;88m-\033[38;2;93;77;83m-\033[38;2;86;70;75m:\033[38;2;64;54;57m:\033[38;2;77;73;74m:\033[38;2;63;63;61m:\033[38;2;62;63;62m:\033[38;2;57;57;58m:\033[38;2;42;42;44m.\033[38;2;38;36;33m.\033[38;2;35;35;37m.\033[38;2;1;1;3m \033[38;2;2;4;3m \033[38;2;6;6;6m \033[38;2;3;1;1m \033[38;2;7;9;8m \033[38;2;8;8;8m \033[38;2;5;5;5m \033[38;2;2;2;2m \033[38;2;2;1;2m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;4m \033[38;2;0;0;2m \033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;0;1m \033[38;2;10;4;6m \033[38;2;13;2;6m \033[38;2;1;0;2m \033[38;2;1;1;3m \033[38;2;2;2;2m \033[38;2;5;5;5m \033[38;2;31;31;31m.\033[38;2;69;60;74m:\033[38;2;60;56;71m:\033[38;2;131;131;141m+\033[38;2;206;206;207m#\033[38;2;252;252;252m@\033[38;2;253;254;255m@\033[38;2;254;254;251m@\033[38;2;254;254;248m@\033[38;2;255;253;254m@\033[38;2;248;246;247m@\033[38;2;252;250;251m@\033[38;2;252;247;249m@\033[38;2;251;249;250m@\033[38;2;249;243;245m@\033[38;2;251;244;246m@\033[38;2;252;245;247m@\033[38;2;253;245;247m@\033[38;2;253;247;247m@\033[38;2;251;245;239m@\033[38;2;251;244;240m@\033[38;2;251;244;237m@\033[38;2;250;243;232m@\033[38;2;249;242;231m@\033[38;2;250;246;238m@\033[38;2;252;247;239m@\033[38;2;251;246;237m@\033[38;2;254;246;240m@\033[38;2;252;242;241m@\033[38;2;253;241;241m@\033[38;2;251;239;239m@\033[38;2;255;243;243m@\033[38;2;255;244;242m@\033[38;2;255;244;242m@\033[38;2;250;241;238m@\033[38;2;253;243;241m@\033[38;2;253;245;240m@\033[38;2;253;242;239m@\033[38;2;253;242;237m@\033[38;2;252;243;238m@\033[38;2;254;246;241m@\033[38;2;254;245;241m@\033[38;2;254;247;239m@\033[38;2;254;245;239m@\033[38;2;249;241;235m@\033[38;2;251;245;241m@\033[38;2;250;244;241m@\033[38;2;252;249;239m@\033[38;2;253;247;238m@\033[38;2;251;245;236m@\033[38;2;250;248;240m@\033[38;2;253;251;241m@\033[38;2;255;251;246m@\033[38;2;255;250;246m@\033[38;2;255;250;249m@\033[38;2;254;248;248m@\033[38;2;255;248;246m@\033[38;2;246;241;238m@\033[38;2;250;246;243m@\033[38;2;252;248;245m@\033[38;2;251;248;247m@\033[38;2;255;253;251m@\033[38;2;253;251;248m@\033[38;2;254;253;247m@\033[38;2;252;251;247m@\033[38;2;255;255;253m@\033[38;2;253;252;250m@\033[38;2;255;255;253m@\033[38;2;253;254;252m@\033[38;2;254;255;252m@\033[38;2;253;255;252m@\033[38;2;254;254;252m@\033[38;2;254;254;252m@\033[38;2;255;252;255m@\033[38;2;255;253;255m@\033[38;2;255;253;251m@\033[38;2;254;253;254m@\033[38;2;252;252;251m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;233;230;231m&\033[38;2;207;202;204m#\033[38;2;174;167;169m*\033[38;2;134;116;120m=\033[38;2;111;91;96m-\033[38;2;73;53;58m:\033[38;2;70;54;59m:\033[38;2;81;71;75m:\033[38;2;74;71;73m:\033[38;2;50;48;49m.\033[38;2;11;9;10m \033[38;2;22;18;19m \033[38;2;1;0;0m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;2m \033[38;2;0;0;4m \033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;0;2m \033[38;2;1;0;2m \033[38;2;1;1;3m \033[38;2;1;1;1m \033[38;2;16;16;16m \033[38;2;56;56;56m:\033[38;2;53;50;68m:\033[38;2;190;187;198m#\033[38;2;251;250;253m@\033[38;2;255;255;253m@\033[38;2;255;255;251m@\033[38;2;253;253;251m@\033[38;2;253;254;249m@\033[38;2;254;254;250m@\033[38;2;253;252;251m@\033[38;2;253;252;248m@\033[38;2;251;252;254m@\033[38;2;254;255;255m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;254;254;254m@\033[38;2;253;255;254m@\033[38;2;252;251;251m@\033[38;2;253;254;253m@\033[38;2;252;250;251m@\033[38;2;254;246;247m@\033[38;2;252;244;236m@\033[38;2;254;244;239m@\033[38;2;252;242;239m@\033[38;2;254;242;241m@\033[38;2;252;242;240m@\033[38;2;253;243;241m@\033[38;2;250;240;238m@\033[38;2;251;241;239m@\033[38;2;250;239;235m@\033[38;2;252;239;233m@\033[38;2;249;238;232m@\033[38;2;252;236;229m@\033[38;2;255;239;232m@\033[38;2;255;241;236m@\033[38;2;251;234;227m@\033[38;2;254;237;229m@\033[38;2;254;237;229m@\033[38;2;250;237;225m@\033[38;2;253;241;227m@\033[38;2;252;242;230m@\033[38;2;255;245;230m@\033[38;2;255;242;222m@\033[38;2;253;240;223m@\033[38;2;253;240;223m@\033[38;2;251;238;221m@\033[38;2;253;240;222m@\033[38;2;254;241;224m@\033[38;2;252;239;230m@\033[38;2;252;239;230m@\033[38;2;252;236;228m@\033[38;2;255;238;229m@\033[38;2;253;236;228m@\033[38;2;250;235;228m@\033[38;2;249;235;226m@\033[38;2;253;240;229m@\033[38;2;254;237;229m@\033[38;2;250;233;225m@\033[38;2;255;238;230m@\033[38;2;254;239;231m@\033[38;2;254;237;229m@\033[38;2;255;241;232m@\033[38;2;255;240;232m@\033[38;2;255;237;230m@\033[38;2;254;238;225m@\033[38;2;252;240;226m@\033[38;2;249;235;226m@\033[38;2;246;232;220m@\033[38;2;251;237;223m@\033[38;2;254;243;230m@\033[38;2;252;242;230m@\033[38;2;247;237;229m@\033[38;2;242;232;223m@\033[38;2;255;248;238m@\033[38;2;252;245;236m@\033[38;2;253;250;245m@\033[38;2;251;253;243m@\033[38;2;252;252;251m@\033[38;2;255;253;255m@\033[38;2;254;255;255m@\033[38;2;253;253;252m@\033[38;2;253;253;255m@\033[38;2;250;253;254m@\033[38;2;252;251;252m@\033[38;2;254;252;253m@\033[38;2;253;252;250m@\033[38;2;251;251;249m@\033[38;2;252;254;251m@\033[38;2;250;255;251m@\033[38;2;251;255;254m@\033[38;2;253;253;254m@\033[38;2;220;215;219m&\033[38;2;152;146;150m+\033[38;2;59;56;58m:\033[38;2;49;47;48m.\033[38;2;25;23;24m \033[38;2;5;3;4m \033[38;2;0;0;2m \033[38;2;1;1;3m \033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;3m \033[38;2;1;0;5m \033[38;2;16;15;21m \033[38;2;62;60;71m:\033[38;2;44;41;60m.\033[38;2;239;238;245m@\033[38;2;251;251;251m@\033[38;2;248;247;252m@\033[38;2;244;244;253m@\033[38;2;244;244;252m@\033[38;2;246;247;252m@\033[38;2;254;254;255m@\033[38;2;145;143;155m+\033[38;2;103;102;109m-\033[38;2;70;70;70m:\033[38;2;74;72;83m:\033[38;2;93;86;94m-\033[38;2;31;24;32m.\033[38;2;94;88;92m-\033[38;2;30;24;28m.\033[38;2;69;63;67m:\033[38;2;75;69;72m:\033[38;2;95;84;88m-\033[38;2;48;33;36m.\033[38;2;165;151;154m*\033[38;2;240;229;231m&\033[38;2;250;248;249m@\033[38;2;252;254;253m@\033[38;2;251;249;249m@\033[38;2;250;245;242m@\033[38;2;249;241;239m@\033[38;2;251;241;239m@\033[38;2;254;243;241m@\033[38;2;252;241;239m@\033[38;2;255;244;242m@\033[38;2;250;240;238m@\033[38;2;249;239;237m@\033[38;2;249;241;236m@\033[38;2;248;239;232m@\033[38;2;251;239;232m@\033[38;2;252;239;231m@\033[38;2;255;239;232m@\033[38;2;255;240;233m@\033[38;2;252;234;227m@\033[38;2;254;238;222m@\033[38;2;255;236;221m@\033[38;2;255;240;224m@\033[38;2;255;240;224m@\033[38;2;255;239;223m@\033[38;2;255;240;224m@\033[38;2;255;238;222m@\033[38;2;251;232;217m@\033[38;2;250;231;215m@\033[38;2;252;233;216m@\033[38;2;254;237;221m@\033[38;2;254;238;223m@\033[38;2;254;237;224m@\033[38;2;255;239;224m@\033[38;2;255;236;221m@\033[38;2;254;238;222m@\033[38;2;255;243;227m@\033[38;2;255;237;223m@\033[38;2;252;239;222m@\033[38;2;255;242;226m@\033[38;2;255;247;230m@\033[38;2;254;243;225m@\033[38;2;244;229;213m&\033[38;2;249;232;214m@\033[38;2;255;239;221m@\033[38;2;249;232;215m@\033[38;2;254;238;222m@\033[38;2;255;247;228m@\033[38;2;254;247;236m@\033[38;2;242;237;225m@\033[38;2;239;236;225m@\033[38;2;250;246;237m@\033[38;2;254;251;246m@\033[38;2;255;253;246m@\033[38;2;253;250;243m@\033[38;2;253;250;243m@\033[38;2;253;253;251m@\033[38;2;251;251;242m@\033[38;2;188;185;148m#\033[38;2;91;87;50m-\033[38;2;41;36;14m.\033[38;2;43;33;7m.\033[38;2;42;33;3m.\033[38;2;121;114;87m=\033[38;2;247;237;226m@\033[38;2;254;243;239m@\033[38;2;253;243;241m@\033[38;2;254;242;242m@\033[38;2;251;235;235m@\033[38;2;251;235;231m@\033[38;2;248;234;233m@\033[38;2;237;231;227m&\033[38;2;253;251;251m@\033[38;2;252;248;247m@\033[38;2;253;253;253m@\033[38;2;253;253;253m@\033[38;2;253;253;253m@\033[38;2;49;49;49m.\033[38;2;47;47;47m.\033[38;2;12;12;14m \033[38;2;1;1;3m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;6;6;6m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;133;133;133m+\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;222;222;222m&\033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;252;252;252m@\033[38;2;48;48;48m.\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;14;14;14m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;251;251;251m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;242;242;242m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;221;221;221m&\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;11;11;11m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;6;6;6m \033[38;2;10;10;10m \033[38;2;4;4;4m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;12;12;12m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;12;12;12m \033[38;2;252;252;252m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;249;249;249m@\033[38;2;254;254;254m@\033[38;2;15;15;15m \033[38;2;7;7;7m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;163;163;163m*\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;122;122;122m=\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;216;216;216m&\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;248;248;248m@\033[38;2;31;31;31m.\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;145;145;145m+\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;249;249;249m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;8;8;8m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;246;246;246m@\033[38;2;248;248;248m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;83;83;83m-\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;245;245;245m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;4;4;4m \033[38;2;253;253;253m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;250;250;250m@\033[38;2;247;247;247m@\033[38;2;4;4;4m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;53;53;53m:\033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;22;22;22m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;27;27;27m.\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;246;246;246m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;5;5;5m \033[38;2;17;17;17m \033[38;2;248;248;248m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;246;246;246m@\033[38;2;24;24;24m \033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;136;136;136m+\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;7;7;7m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;11;11;11m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;11;11;11m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;248;248;248m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;101;101;101m-\033[38;2;5;5;5m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;32;32;32m.\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;11;11;11m \033[38;2;3;3;3m \033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;5;5;5m \033[38;2;248;248;248m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;245;245;245m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;5;5;5m \033[38;2;6;6;6m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;20;20;20m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;1;1;1m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;241;241;241m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;205;205;205m#\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;6;6;6m \033[38;2;2;2;2m \033[38;2;200;200;200m#\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;129;129;129m=\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;5;5;5m \033[38;2;9;9;9m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;46;46;46m.\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;5;5;5m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;7;7;7m \033[38;2;6;6;6m \033[38;2;3;3;3m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;5;5;5m \033[38;2;7;7;7m \033[38;2;18;18;18m \033[38;2;29;29;29m.\033[38;2;38;38;38m.\033[38;2;155;155;155m+\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;249;249;249m@\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;252;252;252m@\033[38;2;249;249;249m@\033[38;2;40;40;40m.\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;250;250;250m@\033[38;2;224;224;224m&\033[38;2;17;17;17m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;143;143;143m+\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;222;222;222m&\033[38;2;6;6;6m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;1;1;1m \033[38;2;246;246;246m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;89;89;89m-\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;251;251;251m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;253;253;253m@\033[38;2;253;253;253m@\033[38;2;225;225;225m&\033[38;2;4;4;4m \033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;11;11;11m \033[38;2;249;249;249m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;252;252;252m@\033[38;2;166;166;166m*\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;135;135;135m+\033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;166;166;166m*\033[38;2;246;246;246m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;246;246;246m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;9;9;9m \033[38;2;250;250;250m@\033[38;2;251;251;251m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;5;5;5m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;9;9;9m \033[38;2;242;242;242m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;249;249;249m@\033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;7;7;7m \033[38;2;12;12;12m \033[38;2;251;251;251m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;217;217;217m&\033[38;2;9;9;9m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;251;251;251m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;250;250;250m@\033[38;2;124;124;124m=\033[38;2;6;6;6m \033[38;2;2;2;2m \033[38;2;3;3;3m \033[38;2;5;5;5m \033[38;2;6;6;6m \033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;221;221;221m&\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;12;12;12m \033[38;2;253;253;253m@\033[38;2;251;251;251m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;11;11;11m \033[38;2;32;32;32m.\033[38;2;250;250;250m@\033[38;2;251;251;251m@\033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;2;2;2m \033[38;2;247;247;247m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;190;190;190m#\033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;201;201;201m#\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;186;186;186m#\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;6;6;6m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;11;11;11m \033[38;2;80;80;80m-\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;80;80;80m-\033[38;2;80;80;80m-\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;3;3;3m \033[38;2;8;8;8m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;53;53;53m:\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;49;49;49m.\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;77;77;77m:\033[38;2;59;59;59m:\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;23;23;23m \033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;7;7;7m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;1;1;1m \033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;250;250;250m@\033[38;2;251;251;251m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;250;250;250m@\033[38;2;20;20;20m \033[38;2;5;5;5m \033[38;2;4;4;4m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;241;241;241m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;162;162;162m*\033[38;2;6;6;6m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;5;5;5m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;11;11;11m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;8;8;8m \033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;64;64;64m:\033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;85;85;85m-\033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;152;152;152m+\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;161;161;161m*\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;50;50;50m.\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;70;70;70m:\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;209;209;209m&\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;2;2;2m \033[38;2;193;193;193m#\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;253;253;253m@\033[38;2;252;252;252m@\033[38;2;252;252;252m@\033[38;2;251;251;251m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;248;248;248m@\033[38;2;88;88;88m-\033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;49;49;49m.\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;244;244;244m@\033[38;2;252;252;252m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;131;131;131m+\033[38;2;253;253;253m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;8;8;8m \033[38;2;247;247;247m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;252;252;252m@\033[38;2;18;18;18m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;6;6;6m \033[38;2;254;254;254m@\033[38;2;250;250;250m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;252;252;252m@\033[38;2;3;3;3m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;4;4;4m \033[38;2;248;248;248m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;251;251;251m@\033[38;2;147;147;147m+\033[38;2;5;5;5m \033[38;2;244;244;244m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;238;238;238m@\033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;199;199;199m#\033[38;2;251;251;251m@\033[38;2;254;254;254m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;253;253;253m@\033[38;2;254;254;254m@\033[38;2;252;252;252m@\033[38;2;253;253;253m@\033[38;2;242;242;242m@\033[38;2;9;9;9m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;4;4;4m \033[38;2;237;237;237m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;254;254;254m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;251;251;251m@\033[38;2;227;227;227m&\033[38;2;0;0;0m \033[38;2;6;6;6m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;3;3;3m \033[38;2;2;2;2m \033[38;2;2;2;2m \033[38;2;4;4;4m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;7;7;7m \033[38;2;17;17;17m \033[38;2;51;51;51m.\033[38;2;70;70;70m:\033[38;2;60;60;60m:\033[38;2;38;38;38m.\033[38;2;8;8;8m \033[38;2;4;4;4m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;1;1;1m \033[38;2;2;2;2m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;3;3;3m \033[38;2;5;5;5m \033[38;2;27;27;27m.\033[38;2;54;54;54m:\033[38;2;74;74;74m:\033[38;2;58;58;58m:\033[38;2;20;20;20m \033[38;2;5;5;5m \033[38;2;1;1;1m \033[38;2;1;1;1m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
        $display("\033[38;2;0;0;2m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[38;2;0;0;0m \033[0m");
    end
    endtask

endmodule
